`timescale 1ns/100ps

module data_rom ( 
// write input and output here.
input           clk;
input           rst_n;
input           ena;
);
always @(posedge clk) begin 
    case(address)
        'd0 :data = 'd1;
        'd1 :data = 'd0;
        'd2 :data = 'd0;
        'd3 :data = 'd0;
        'd4 :data = 'd1;
        'd5 :data = 'd1;
        'd6 :data = 'd1;
        'd7 :data = 'd1;
        'd8 :data = 'd1;
        'd9 :data = 'd1;
        'd10 :data = 'd1;
        'd11 :data = 'd1;
        'd12 :data = 'd0;
        'd13 :data = 'd0;
        'd14 :data = 'd0;
        'd15 :data = 'd1;
        'd16 :data = 'd1;
        'd17 :data = 'd1;
        'd18 :data = 'd1;
        'd19 :data = 'd1;
        'd20 :data = 'd1;
        'd21 :data = 'd1;
        'd22 :data = 'd0;
        'd23 :data = 'd0;
        'd24 :data = 'd0;
        'd25 :data = 'd1;
        'd26 :data = 'd1;
        'd27 :data = 'd1;
        'd28 :data = 'd1;
        'd29 :data = 'd0;
        'd30 :data = 'd0;
        'd31 :data = 'd1;
        'd32 :data = 'd1;
        'd33 :data = 'd0;
        'd34 :data = 'd0;
        'd35 :data = 'd1;
        'd36 :data = 'd1;
        'd37 :data = 'd0;
        'd38 :data = 'd1;
        'd39 :data = 'd1;
        'd40 :data = 'd1;
        'd41 :data = 'd1;
        'd42 :data = 'd1;
        'd43 :data = 'd0;
        'd44 :data = 'd0;
        'd45 :data = 'd0;
        'd46 :data = 'd0;
        'd47 :data = 'd0;
        'd48 :data = 'd1;
        'd49 :data = 'd0;
        'd50 :data = 'd1;
        'd51 :data = 'd0;
        'd52 :data = 'd1;
        'd53 :data = 'd1;
        'd54 :data = 'd1;
        'd55 :data = 'd0;
        'd56 :data = 'd0;
        'd57 :data = 'd0;
        'd58 :data = 'd1;
        'd59 :data = 'd1;
        'd60 :data = 'd0;
        'd61 :data = 'd0;
        'd62 :data = 'd1;
        'd63 :data = 'd0;
        'd64 :data = 'd0;
        'd65 :data = 'd1;
        'd66 :data = 'd1;
        'd67 :data = 'd1;
        'd68 :data = 'd1;
        'd69 :data = 'd1;
        'd70 :data = 'd1;
        'd71 :data = 'd0;
        'd72 :data = 'd0;
        'd73 :data = 'd1;
        'd74 :data = 'd1;
        'd75 :data = 'd0;
        'd76 :data = 'd0;
        'd77 :data = 'd1;
        'd78 :data = 'd0;
        'd79 :data = 'd1;
        'd80 :data = 'd1;
        'd81 :data = 'd1;
        'd82 :data = 'd0;
        'd83 :data = 'd1;
        'd84 :data = 'd0;
        'd85 :data = 'd0;
        'd86 :data = 'd0;
        'd87 :data = 'd0;
        'd88 :data = 'd1;
        'd89 :data = 'd0;
        'd90 :data = 'd1;
        'd91 :data = 'd1;
        'd92 :data = 'd1;
        'd93 :data = 'd1;
        'd94 :data = 'd0;
        'd95 :data = 'd1;
        'd96 :data = 'd0;
        'd97 :data = 'd1;
        'd98 :data = 'd1;
        'd99 :data = 'd0;
        'd100 :data = 'd0;
        'd101 :data = 'd0;
        'd102 :data = 'd1;
        'd103 :data = 'd0;
        'd104 :data = 'd0;
        'd105 :data = 'd1;
        'd106 :data = 'd1;
        'd107 :data = 'd1;
        'd108 :data = 'd1;
        'd109 :data = 'd1;
        'd110 :data = 'd1;
        'd111 :data = 'd0;
        'd112 :data = 'd1;
        'd113 :data = 'd0;
        'd114 :data = 'd0;
        'd115 :data = 'd1;
        'd116 :data = 'd1;
        'd117 :data = 'd1;
        'd118 :data = 'd1;
        'd119 :data = 'd0;
        'd120 :data = 'd1;
        'd121 :data = 'd1;
        'd122 :data = 'd0;
        'd123 :data = 'd1;
        'd124 :data = 'd1;
        'd125 :data = 'd1;
        'd126 :data = 'd0;
        'd127 :data = 'd0;
        'd128 :data = 'd0;
        'd129 :data = 'd0;
        'd130 :data = 'd0;
        'd131 :data = 'd0;
        'd132 :data = 'd1;
        'd133 :data = 'd1;
        'd134 :data = 'd1;
        'd135 :data = 'd0;
        'd136 :data = 'd0;
        'd137 :data = 'd1;
        'd138 :data = 'd1;
        'd139 :data = 'd0;
        'd140 :data = 'd0;
        'd141 :data = 'd1;
        'd142 :data = 'd0;
        'd143 :data = 'd0;
        'd144 :data = 'd0;
        'd145 :data = 'd1;
        'd146 :data = 'd0;
        'd147 :data = 'd1;
        'd148 :data = 'd0;
        'd149 :data = 'd0;
        'd150 :data = 'd1;
        'd151 :data = 'd1;
        'd152 :data = 'd0;
        'd153 :data = 'd0;
        'd154 :data = 'd0;
        'd155 :data = 'd1;
        'd156 :data = 'd1;
        'd157 :data = 'd1;
        'd158 :data = 'd0;
        'd159 :data = 'd1;
        'd160 :data = 'd0;
        'd161 :data = 'd0;
        'd162 :data = 'd0;
        'd163 :data = 'd0;
        'd164 :data = 'd1;
        'd165 :data = 'd1;
        'd166 :data = 'd1;
        'd167 :data = 'd1;
        'd168 :data = 'd0;
        'd169 :data = 'd1;
        'd170 :data = 'd1;
        'd171 :data = 'd0;
        'd172 :data = 'd1;
        'd173 :data = 'd1;
        'd174 :data = 'd1;
        'd175 :data = 'd0;
        'd176 :data = 'd1;
        'd177 :data = 'd1;
        'd178 :data = 'd1;
        'd179 :data = 'd0;
        'd180 :data = 'd0;
        'd181 :data = 'd0;
        'd182 :data = 'd1;
        'd183 :data = 'd0;
        'd184 :data = 'd0;
        'd185 :data = 'd1;
        'd186 :data = 'd0;
        'd187 :data = 'd1;
        'd188 :data = 'd0;
        'd189 :data = 'd0;
        'd190 :data = 'd1;
        'd191 :data = 'd1;
        'd192 :data = 'd0;
        'd193 :data = 'd0;
        'd194 :data = 'd1;
        'd195 :data = 'd0;
        'd196 :data = 'd0;
        'd197 :data = 'd0;
        'd198 :data = 'd0;
        'd199 :data = 'd1;
        'd200 :data = 'd1;
        'd201 :data = 'd0;
        'd202 :data = 'd0;
        'd203 :data = 'd1;
        'd204 :data = 'd0;
        'd205 :data = 'd0;
        'd206 :data = 'd1;
        'd207 :data = 'd0;
        'd208 :data = 'd1;
        'd209 :data = 'd0;
        'd210 :data = 'd1;
        'd211 :data = 'd0;
        'd212 :data = 'd1;
        'd213 :data = 'd1;
        'd214 :data = 'd0;
        'd215 :data = 'd1;
        'd216 :data = 'd0;
        'd217 :data = 'd1;
        'd218 :data = 'd0;
        'd219 :data = 'd0;
        'd220 :data = 'd0;
        'd221 :data = 'd0;
        'd222 :data = 'd0;
        'd223 :data = 'd1;
        'd224 :data = 'd0;
        'd225 :data = 'd0;
        'd226 :data = 'd1;
        'd227 :data = 'd0;
        'd228 :data = 'd1;
        'd229 :data = 'd1;
        'd230 :data = 'd0;
        'd231 :data = 'd0;
        'd232 :data = 'd0;
        'd233 :data = 'd0;
        'd234 :data = 'd0;
        'd235 :data = 'd0;
        'd236 :data = 'd0;
        'd237 :data = 'd0;
        'd238 :data = 'd1;
        'd239 :data = 'd1;
        'd240 :data = 'd1;
        'd241 :data = 'd1;
        'd242 :data = 'd0;
        'd243 :data = 'd0;
        'd244 :data = 'd0;
        'd245 :data = 'd1;
        'd246 :data = 'd1;
        'd247 :data = 'd1;
        'd248 :data = 'd0;
        'd249 :data = 'd1;
        'd250 :data = 'd0;
        'd251 :data = 'd1;
        'd252 :data = 'd1;
        'd253 :data = 'd1;
        'd254 :data = 'd0;
        'd255 :data = 'd0;
        'd256 :data = 'd0;
        'd257 :data = 'd0;
        'd258 :data = 'd0;
        'd259 :data = 'd0;
        'd260 :data = 'd1;
        'd261 :data = 'd1;
        'd262 :data = 'd1;
        'd263 :data = 'd0;
        'd264 :data = 'd1;
        'd265 :data = 'd0;
        'd266 :data = 'd1;
        'd267 :data = 'd0;
        'd268 :data = 'd0;
        'd269 :data = 'd1;
        'd270 :data = 'd1;
        'd271 :data = 'd0;
        'd272 :data = 'd0;
        'd273 :data = 'd1;
        'd274 :data = 'd0;
        'd275 :data = 'd0;
        'd276 :data = 'd1;
        'd277 :data = 'd1;
        'd278 :data = 'd1;
        'd279 :data = 'd0;
        'd280 :data = 'd1;
        'd281 :data = 'd1;
        'd282 :data = 'd1;
        'd283 :data = 'd1;
        'd284 :data = 'd1;
        'd285 :data = 'd0;
        'd286 :data = 'd0;
        'd287 :data = 'd0;
        'd288 :data = 'd0;
        'd289 :data = 'd1;
        'd290 :data = 'd1;
        'd291 :data = 'd0;
        'd292 :data = 'd0;
        'd293 :data = 'd0;
        'd294 :data = 'd1;
        'd295 :data = 'd0;
        'd296 :data = 'd1;
        'd297 :data = 'd1;
        'd298 :data = 'd0;
        'd299 :data = 'd0;
        'd300 :data = 'd0;
        'd301 :data = 'd1;
        'd302 :data = 'd0;
        'd303 :data = 'd1;
        'd304 :data = 'd0;
        'd305 :data = 'd1;
        'd306 :data = 'd0;
        'd307 :data = 'd1;
        'd308 :data = 'd1;
        'd309 :data = 'd0;
        'd310 :data = 'd0;
        'd311 :data = 'd1;
        'd312 :data = 'd1;
        'd313 :data = 'd0;
        'd314 :data = 'd0;
        'd315 :data = 'd0;
        'd316 :data = 'd1;
        'd317 :data = 'd0;
        'd318 :data = 'd0;
        'd319 :data = 'd1;
        'd320 :data = 'd0;
        'd321 :data = 'd0;
        'd322 :data = 'd1;
        'd323 :data = 'd0;
        'd324 :data = 'd1;
        'd325 :data = 'd0;
        'd326 :data = 'd1;
        'd327 :data = 'd0;
        'd328 :data = 'd0;
        'd329 :data = 'd0;
        'd330 :data = 'd1;
        'd331 :data = 'd0;
        'd332 :data = 'd1;
        'd333 :data = 'd0;
        'd334 :data = 'd0;
        'd335 :data = 'd1;
        'd336 :data = 'd1;
        'd337 :data = 'd0;
        'd338 :data = 'd0;
        'd339 :data = 'd1;
        'd340 :data = 'd0;
        'd341 :data = 'd0;
        'd342 :data = 'd0;
        'd343 :data = 'd0;
        'd344 :data = 'd0;
        'd345 :data = 'd0;
        'd346 :data = 'd0;
        'd347 :data = 'd0;
        'd348 :data = 'd0;
        'd349 :data = 'd1;
        'd350 :data = 'd0;
        'd351 :data = 'd1;
        'd352 :data = 'd0;
        'd353 :data = 'd1;
        'd354 :data = 'd1;
        'd355 :data = 'd0;
        'd356 :data = 'd1;
        'd357 :data = 'd0;
        'd358 :data = 'd1;
        'd359 :data = 'd0;
        'd360 :data = 'd1;
        'd361 :data = 'd0;
        'd362 :data = 'd0;
        'd363 :data = 'd1;
        'd364 :data = 'd1;
        'd365 :data = 'd1;
        'd366 :data = 'd1;
        'd367 :data = 'd0;
        'd368 :data = 'd0;
        'd369 :data = 'd1;
        'd370 :data = 'd1;
        'd371 :data = 'd0;
        'd372 :data = 'd0;
        'd373 :data = 'd0;
        'd374 :data = 'd1;
        'd375 :data = 'd1;
        'd376 :data = 'd0;
        'd377 :data = 'd1;
        'd378 :data = 'd0;
        'd379 :data = 'd0;
        'd380 :data = 'd1;
        'd381 :data = 'd1;
        'd382 :data = 'd1;
        'd383 :data = 'd0;
        'd384 :data = 'd1;
        'd385 :data = 'd1;
        'd386 :data = 'd0;
        'd387 :data = 'd1;
        'd388 :data = 'd0;
        'd389 :data = 'd1;
        'd390 :data = 'd1;
        'd391 :data = 'd1;
        'd392 :data = 'd1;
        'd393 :data = 'd0;
        'd394 :data = 'd0;
        'd395 :data = 'd1;
        'd396 :data = 'd1;
        'd397 :data = 'd0;
        'd398 :data = 'd0;
        'd399 :data = 'd1;
        'd400 :data = 'd1;
        'd401 :data = 'd0;
        'd402 :data = 'd0;
        'd403 :data = 'd0;
        'd404 :data = 'd0;
        'd405 :data = 'd1;
        'd406 :data = 'd1;
        'd407 :data = 'd0;
        'd408 :data = 'd0;
        'd409 :data = 'd0;
        'd410 :data = 'd0;
        'd411 :data = 'd1;
        'd412 :data = 'd1;
        'd413 :data = 'd1;
        'd414 :data = 'd1;
        'd415 :data = 'd1;
        'd416 :data = 'd0;
        'd417 :data = 'd1;
        'd418 :data = 'd1;
        'd419 :data = 'd0;
        'd420 :data = 'd1;
        'd421 :data = 'd1;
        'd422 :data = 'd1;
        'd423 :data = 'd1;
        'd424 :data = 'd0;
        'd425 :data = 'd1;
        'd426 :data = 'd0;
        'd427 :data = 'd0;
        'd428 :data = 'd0;
        'd429 :data = 'd0;
        'd430 :data = 'd1;
        'd431 :data = 'd1;
        'd432 :data = 'd1;
        'd433 :data = 'd1;
        'd434 :data = 'd1;
        'd435 :data = 'd0;
        'd436 :data = 'd0;
        'd437 :data = 'd0;
        'd438 :data = 'd0;
        'd439 :data = 'd1;
        'd440 :data = 'd1;
        'd441 :data = 'd0;
        'd442 :data = 'd1;
        'd443 :data = 'd1;
        'd444 :data = 'd0;
        'd445 :data = 'd1;
        'd446 :data = 'd0;
        'd447 :data = 'd0;
        'd448 :data = 'd1;
        'd449 :data = 'd0;
        'd450 :data = 'd0;
        'd451 :data = 'd0;
        'd452 :data = 'd0;
        'd453 :data = 'd1;
        'd454 :data = 'd0;
        'd455 :data = 'd0;
        'd456 :data = 'd1;
        'd457 :data = 'd1;
        'd458 :data = 'd0;
        'd459 :data = 'd1;
        'd460 :data = 'd1;
        'd461 :data = 'd0;
        'd462 :data = 'd1;
        'd463 :data = 'd0;
        'd464 :data = 'd1;
        'd465 :data = 'd0;
        'd466 :data = 'd0;
        'd467 :data = 'd1;
        'd468 :data = 'd0;
        'd469 :data = 'd0;
        'd470 :data = 'd1;
        'd471 :data = 'd1;
        'd472 :data = 'd1;
        'd473 :data = 'd0;
        'd474 :data = 'd0;
        'd475 :data = 'd1;
        'd476 :data = 'd1;
        'd477 :data = 'd0;
        'd478 :data = 'd1;
        'd479 :data = 'd1;
        'd480 :data = 'd1;
        'd481 :data = 'd0;
        'd482 :data = 'd1;
        'd483 :data = 'd0;
        'd484 :data = 'd1;
        'd485 :data = 'd0;
        'd486 :data = 'd1;
        'd487 :data = 'd0;
        'd488 :data = 'd1;
        'd489 :data = 'd1;
        'd490 :data = 'd0;
        'd491 :data = 'd1;
        'd492 :data = 'd1;
        'd493 :data = 'd1;
        'd494 :data = 'd1;
        'd495 :data = 'd1;
        'd496 :data = 'd1;
        'd497 :data = 'd1;
        'd498 :data = 'd0;
        'd499 :data = 'd1;
        'd500 :data = 'd0;
        'd501 :data = 'd0;
        'd502 :data = 'd1;
        'd503 :data = 'd1;
        'd504 :data = 'd0;
        'd505 :data = 'd0;
        'd506 :data = 'd0;
        'd507 :data = 'd0;
        'd508 :data = 'd1;
        'd509 :data = 'd0;
        'd510 :data = 'd0;
        'd511 :data = 'd0;
        'd512 :data = 'd0;
        'd513 :data = 'd0;
        'd514 :data = 'd1;
        'd515 :data = 'd0;
        'd516 :data = 'd1;
        'd517 :data = 'd1;
        'd518 :data = 'd1;
        'd519 :data = 'd1;
        'd520 :data = 'd0;
        'd521 :data = 'd0;
        'd522 :data = 'd1;
        'd523 :data = 'd1;
        'd524 :data = 'd1;
        'd525 :data = 'd0;
        'd526 :data = 'd0;
        'd527 :data = 'd0;
        'd528 :data = 'd1;
        'd529 :data = 'd1;
        'd530 :data = 'd1;
        'd531 :data = 'd0;
        'd532 :data = 'd1;
        'd533 :data = 'd1;
        'd534 :data = 'd1;
        'd535 :data = 'd0;
        'd536 :data = 'd1;
        'd537 :data = 'd0;
        'd538 :data = 'd0;
        'd539 :data = 'd1;
        'd540 :data = 'd1;
        'd541 :data = 'd1;
        'd542 :data = 'd0;
        'd543 :data = 'd0;
        'd544 :data = 'd0;
        'd545 :data = 'd0;
        'd546 :data = 'd1;
        'd547 :data = 'd1;
        'd548 :data = 'd1;
        'd549 :data = 'd0;
        'd550 :data = 'd0;
        'd551 :data = 'd0;
        'd552 :data = 'd0;
        'd553 :data = 'd1;
        'd554 :data = 'd1;
        'd555 :data = 'd0;
        'd556 :data = 'd1;
        'd557 :data = 'd0;
        'd558 :data = 'd0;
        'd559 :data = 'd1;
        'd560 :data = 'd0;
        'd561 :data = 'd0;
        'd562 :data = 'd0;
        'd563 :data = 'd1;
        'd564 :data = 'd0;
        'd565 :data = 'd1;
        'd566 :data = 'd0;
        'd567 :data = 'd1;
        'd568 :data = 'd1;
        'd569 :data = 'd0;
        'd570 :data = 'd1;
        'd571 :data = 'd0;
        'd572 :data = 'd1;
        'd573 :data = 'd1;
        'd574 :data = 'd0;
        'd575 :data = 'd1;
        'd576 :data = 'd1;
        'd577 :data = 'd0;
        'd578 :data = 'd1;
        'd579 :data = 'd0;
        'd580 :data = 'd0;
        'd581 :data = 'd0;
        'd582 :data = 'd1;
        'd583 :data = 'd0;
        'd584 :data = 'd1;
        'd585 :data = 'd1;
        'd586 :data = 'd1;
        'd587 :data = 'd0;
        'd588 :data = 'd0;
        'd589 :data = 'd1;
        'd590 :data = 'd1;
        'd591 :data = 'd0;
        'd592 :data = 'd0;
        'd593 :data = 'd1;
        'd594 :data = 'd1;
        'd595 :data = 'd0;
        'd596 :data = 'd1;
        'd597 :data = 'd0;
        'd598 :data = 'd1;
        'd599 :data = 'd0;
        'd600 :data = 'd0;
        'd601 :data = 'd1;
        'd602 :data = 'd1;
        'd603 :data = 'd0;
        'd604 :data = 'd1;
        'd605 :data = 'd1;
        'd606 :data = 'd1;
        'd607 :data = 'd1;
        'd608 :data = 'd0;
        'd609 :data = 'd0;
        'd610 :data = 'd1;
        'd611 :data = 'd0;
        'd612 :data = 'd0;
        'd613 :data = 'd1;
        'd614 :data = 'd1;
        'd615 :data = 'd0;
        'd616 :data = 'd1;
        'd617 :data = 'd0;
        'd618 :data = 'd0;
        'd619 :data = 'd1;
        'd620 :data = 'd0;
        'd621 :data = 'd0;
        'd622 :data = 'd1;
        'd623 :data = 'd1;
        'd624 :data = 'd1;
        'd625 :data = 'd0;
        'd626 :data = 'd1;
        'd627 :data = 'd1;
        'd628 :data = 'd1;
        'd629 :data = 'd1;
        'd630 :data = 'd1;
        'd631 :data = 'd1;
        'd632 :data = 'd0;
        'd633 :data = 'd0;
        'd634 :data = 'd1;
        'd635 :data = 'd1;
        'd636 :data = 'd0;
        'd637 :data = 'd1;
        'd638 :data = 'd1;
        'd639 :data = 'd1;
        'd640 :data = 'd0;
        'd641 :data = 'd0;
        'd642 :data = 'd0;
        'd643 :data = 'd1;
        'd644 :data = 'd1;
        'd645 :data = 'd0;
        'd646 :data = 'd1;
        'd647 :data = 'd1;
        'd648 :data = 'd0;
        'd649 :data = 'd1;
        'd650 :data = 'd0;
        'd651 :data = 'd0;
        'd652 :data = 'd0;
        'd653 :data = 'd0;
        'd654 :data = 'd0;
        'd655 :data = 'd0;
        'd656 :data = 'd1;
        'd657 :data = 'd1;
        'd658 :data = 'd1;
        'd659 :data = 'd1;
        'd660 :data = 'd0;
        'd661 :data = 'd1;
        'd662 :data = 'd0;
        'd663 :data = 'd1;
        'd664 :data = 'd1;
        'd665 :data = 'd0;
        'd666 :data = 'd1;
        'd667 :data = 'd0;
        'd668 :data = 'd0;
        'd669 :data = 'd0;
        'd670 :data = 'd1;
        'd671 :data = 'd0;
        'd672 :data = 'd1;
        'd673 :data = 'd0;
        'd674 :data = 'd1;
        'd675 :data = 'd1;
        'd676 :data = 'd1;
        'd677 :data = 'd0;
        'd678 :data = 'd1;
        'd679 :data = 'd1;
        'd680 :data = 'd0;
        'd681 :data = 'd1;
        'd682 :data = 'd1;
        'd683 :data = 'd1;
        'd684 :data = 'd1;
        'd685 :data = 'd1;
        'd686 :data = 'd1;
        'd687 :data = 'd0;
        'd688 :data = 'd0;
        'd689 :data = 'd0;
        'd690 :data = 'd0;
        'd691 :data = 'd1;
        'd692 :data = 'd0;
        'd693 :data = 'd1;
        'd694 :data = 'd1;
        'd695 :data = 'd1;
        'd696 :data = 'd1;
        'd697 :data = 'd0;
        'd698 :data = 'd0;
        'd699 :data = 'd0;
        'd700 :data = 'd0;
        'd701 :data = 'd1;
        'd702 :data = 'd1;
        'd703 :data = 'd1;
        'd704 :data = 'd0;
        'd705 :data = 'd0;
        'd706 :data = 'd1;
        'd707 :data = 'd1;
        'd708 :data = 'd0;
        'd709 :data = 'd0;
        'd710 :data = 'd0;
        'd711 :data = 'd1;
        'd712 :data = 'd1;
        'd713 :data = 'd1;
        'd714 :data = 'd1;
        'd715 :data = 'd0;
        'd716 :data = 'd1;
        'd717 :data = 'd1;
        'd718 :data = 'd1;
        'd719 :data = 'd1;
        'd720 :data = 'd0;
        'd721 :data = 'd0;
        'd722 :data = 'd0;
        'd723 :data = 'd0;
        'd724 :data = 'd1;
        'd725 :data = 'd0;
        'd726 :data = 'd1;
        'd727 :data = 'd1;
        'd728 :data = 'd0;
        'd729 :data = 'd0;
        'd730 :data = 'd0;
        'd731 :data = 'd1;
        'd732 :data = 'd1;
        'd733 :data = 'd1;
        'd734 :data = 'd0;
        'd735 :data = 'd0;
        'd736 :data = 'd0;
        'd737 :data = 'd1;
        'd738 :data = 'd1;
        'd739 :data = 'd0;
        'd740 :data = 'd1;
        'd741 :data = 'd0;
        'd742 :data = 'd0;
        'd743 :data = 'd1;
        'd744 :data = 'd1;
        'd745 :data = 'd0;
        'd746 :data = 'd0;
        'd747 :data = 'd0;
        'd748 :data = 'd1;
        'd749 :data = 'd0;
        'd750 :data = 'd0;
        'd751 :data = 'd0;
        'd752 :data = 'd0;
        'd753 :data = 'd1;
        'd754 :data = 'd0;
        'd755 :data = 'd0;
        'd756 :data = 'd1;
        'd757 :data = 'd1;
        'd758 :data = 'd0;
        'd759 :data = 'd0;
        'd760 :data = 'd1;
        'd761 :data = 'd0;
        'd762 :data = 'd1;
        'd763 :data = 'd1;
        'd764 :data = 'd1;
        'd765 :data = 'd1;
        'd766 :data = 'd1;
        'd767 :data = 'd0;
        'd768 :data = 'd0;
        'd769 :data = 'd1;
        'd770 :data = 'd1;
        'd771 :data = 'd0;
        'd772 :data = 'd1;
        'd773 :data = 'd0;
        'd774 :data = 'd0;
        'd775 :data = 'd1;
        'd776 :data = 'd1;
        'd777 :data = 'd1;
        'd778 :data = 'd0;
        'd779 :data = 'd0;
        'd780 :data = 'd0;
        'd781 :data = 'd1;
        'd782 :data = 'd0;
        'd783 :data = 'd0;
        'd784 :data = 'd0;
        'd785 :data = 'd0;
        'd786 :data = 'd1;
        'd787 :data = 'd1;
        'd788 :data = 'd1;
        'd789 :data = 'd0;
        'd790 :data = 'd1;
        'd791 :data = 'd1;
        'd792 :data = 'd1;
        'd793 :data = 'd0;
        'd794 :data = 'd0;
        'd795 :data = 'd1;
        'd796 :data = 'd1;
        'd797 :data = 'd0;
        'd798 :data = 'd1;
        'd799 :data = 'd0;
        'd800 :data = 'd0;
        'd801 :data = 'd1;
        'd802 :data = 'd1;
        'd803 :data = 'd0;
        'd804 :data = 'd0;
        'd805 :data = 'd0;
        'd806 :data = 'd1;
        'd807 :data = 'd0;
        'd808 :data = 'd0;
        'd809 :data = 'd1;
        'd810 :data = 'd0;
        'd811 :data = 'd0;
        'd812 :data = 'd1;
        'd813 :data = 'd1;
        'd814 :data = 'd0;
        'd815 :data = 'd1;
        'd816 :data = 'd0;
        'd817 :data = 'd0;
        'd818 :data = 'd0;
        'd819 :data = 'd1;
        'd820 :data = 'd0;
        'd821 :data = 'd0;
        'd822 :data = 'd1;
        'd823 :data = 'd1;
        'd824 :data = 'd0;
        'd825 :data = 'd1;
        'd826 :data = 'd1;
        'd827 :data = 'd0;
        'd828 :data = 'd1;
        'd829 :data = 'd0;
        'd830 :data = 'd0;
        'd831 :data = 'd0;
        'd832 :data = 'd0;
        'd833 :data = 'd0;
        'd834 :data = 'd0;
        'd835 :data = 'd1;
        'd836 :data = 'd0;
        'd837 :data = 'd1;
        'd838 :data = 'd1;
        'd839 :data = 'd1;
        'd840 :data = 'd0;
        'd841 :data = 'd1;
        'd842 :data = 'd0;
        'd843 :data = 'd1;
        'd844 :data = 'd0;
        'd845 :data = 'd1;
        'd846 :data = 'd0;
        'd847 :data = 'd1;
        'd848 :data = 'd1;
        'd849 :data = 'd0;
        'd850 :data = 'd0;
        'd851 :data = 'd0;
        'd852 :data = 'd1;
        'd853 :data = 'd0;
        'd854 :data = 'd1;
        'd855 :data = 'd0;
        'd856 :data = 'd0;
        'd857 :data = 'd1;
        'd858 :data = 'd1;
        'd859 :data = 'd1;
        'd860 :data = 'd0;
        'd861 :data = 'd0;
        'd862 :data = 'd1;
        'd863 :data = 'd1;
        'd864 :data = 'd1;
        'd865 :data = 'd1;
        'd866 :data = 'd0;
        'd867 :data = 'd0;
        'd868 :data = 'd0;
        'd869 :data = 'd1;
        'd870 :data = 'd1;
        'd871 :data = 'd0;
        'd872 :data = 'd0;
        'd873 :data = 'd1;
        'd874 :data = 'd0;
        'd875 :data = 'd1;
        'd876 :data = 'd1;
        'd877 :data = 'd0;
        'd878 :data = 'd1;
        'd879 :data = 'd0;
        'd880 :data = 'd1;
        'd881 :data = 'd0;
        'd882 :data = 'd0;
        'd883 :data = 'd0;
        'd884 :data = 'd1;
        'd885 :data = 'd1;
        'd886 :data = 'd0;
        'd887 :data = 'd1;
        'd888 :data = 'd0;
        'd889 :data = 'd1;
        'd890 :data = 'd1;
        'd891 :data = 'd1;
        'd892 :data = 'd1;
        'd893 :data = 'd0;
        'd894 :data = 'd0;
        'd895 :data = 'd1;
        'd896 :data = 'd1;
        'd897 :data = 'd0;
        'd898 :data = 'd1;
        'd899 :data = 'd0;
        'd900 :data = 'd0;
        'd901 :data = 'd1;
        'd902 :data = 'd0;
        'd903 :data = 'd1;
        'd904 :data = 'd0;
        'd905 :data = 'd1;
        'd906 :data = 'd0;
        'd907 :data = 'd0;
        'd908 :data = 'd0;
        'd909 :data = 'd1;
        'd910 :data = 'd1;
        'd911 :data = 'd0;
        'd912 :data = 'd1;
        'd913 :data = 'd1;
        'd914 :data = 'd0;
        'd915 :data = 'd0;
        'd916 :data = 'd1;
        'd917 :data = 'd0;
        'd918 :data = 'd1;
        'd919 :data = 'd0;
        'd920 :data = 'd1;
        'd921 :data = 'd1;
        'd922 :data = 'd0;
        'd923 :data = 'd1;
        'd924 :data = 'd0;
        'd925 :data = 'd1;
        'd926 :data = 'd1;
        'd927 :data = 'd1;
        'd928 :data = 'd1;
        'd929 :data = 'd1;
        'd930 :data = 'd0;
        'd931 :data = 'd0;
        'd932 :data = 'd0;
        'd933 :data = 'd0;
        'd934 :data = 'd0;
        'd935 :data = 'd1;
        'd936 :data = 'd1;
        'd937 :data = 'd1;
        'd938 :data = 'd0;
        'd939 :data = 'd1;
        'd940 :data = 'd1;
        'd941 :data = 'd1;
        'd942 :data = 'd0;
        'd943 :data = 'd0;
        'd944 :data = 'd0;
        'd945 :data = 'd0;
        'd946 :data = 'd1;
        'd947 :data = 'd1;
        'd948 :data = 'd0;
        'd949 :data = 'd0;
        'd950 :data = 'd0;
        'd951 :data = 'd1;
        'd952 :data = 'd0;
        'd953 :data = 'd1;
        'd954 :data = 'd1;
        'd955 :data = 'd1;
        'd956 :data = 'd1;
        'd957 :data = 'd0;
        'd958 :data = 'd1;
        'd959 :data = 'd1;
        'd960 :data = 'd1;
        'd961 :data = 'd0;
        'd962 :data = 'd0;
        'd963 :data = 'd1;
        'd964 :data = 'd0;
        'd965 :data = 'd1;
        'd966 :data = 'd1;
        'd967 :data = 'd1;
        'd968 :data = 'd0;
        'd969 :data = 'd1;
        'd970 :data = 'd0;
        'd971 :data = 'd0;
        'd972 :data = 'd1;
        'd973 :data = 'd0;
        'd974 :data = 'd0;
        'd975 :data = 'd0;
        'd976 :data = 'd1;
        'd977 :data = 'd1;
        'd978 :data = 'd0;
        'd979 :data = 'd0;
        'd980 :data = 'd0;
        'd981 :data = 'd1;
        'd982 :data = 'd1;
        'd983 :data = 'd1;
        'd984 :data = 'd1;
        'd985 :data = 'd0;
        'd986 :data = 'd0;
        'd987 :data = 'd0;
        'd988 :data = 'd1;
        'd989 :data = 'd0;
        'd990 :data = 'd0;
        'd991 :data = 'd0;
        'd992 :data = 'd0;
        'd993 :data = 'd1;
        'd994 :data = 'd1;
        'd995 :data = 'd0;
        'd996 :data = 'd1;
        'd997 :data = 'd1;
        'd998 :data = 'd0;
        'd999 :data = 'd0;
        'd1000 :data = 'd1;
        'd1001 :data = 'd1;
        'd1002 :data = 'd1;
        'd1003 :data = 'd1;
        'd1004 :data = 'd1;
        'd1005 :data = 'd1;
        'd1006 :data = 'd0;
        'd1007 :data = 'd1;
        'd1008 :data = 'd1;
        'd1009 :data = 'd1;
        'd1010 :data = 'd0;
        'd1011 :data = 'd1;
        'd1012 :data = 'd1;
        'd1013 :data = 'd1;
        'd1014 :data = 'd0;
        'd1015 :data = 'd0;
        'd1016 :data = 'd1;
        'd1017 :data = 'd1;
        'd1018 :data = 'd1;
        'd1019 :data = 'd1;
        'd1020 :data = 'd1;
        'd1021 :data = 'd1;
        'd1022 :data = 'd0;
        'd1023 :data = 'd0;
        'd1024 :data = 'd1;
        'd1025 :data = 'd1;
        'd1026 :data = 'd0;
        'd1027 :data = 'd0;
        'd1028 :data = 'd1;
        'd1029 :data = 'd0;
        'd1030 :data = 'd0;
        'd1031 :data = 'd1;
        'd1032 :data = 'd1;
        'd1033 :data = 'd1;
        'd1034 :data = 'd0;
        'd1035 :data = 'd1;
        'd1036 :data = 'd1;
        'd1037 :data = 'd1;
        'd1038 :data = 'd1;
        'd1039 :data = 'd1;
        'd1040 :data = 'd1;
        'd1041 :data = 'd1;
        'd1042 :data = 'd0;
        'd1043 :data = 'd1;
        'd1044 :data = 'd0;
        'd1045 :data = 'd1;
        'd1046 :data = 'd1;
        'd1047 :data = 'd0;
        'd1048 :data = 'd1;
        'd1049 :data = 'd1;
        'd1050 :data = 'd1;
        'd1051 :data = 'd1;
        'd1052 :data = 'd0;
        'd1053 :data = 'd0;
        'd1054 :data = 'd1;
        'd1055 :data = 'd1;
        'd1056 :data = 'd1;
        'd1057 :data = 'd1;
        'd1058 :data = 'd0;
        'd1059 :data = 'd1;
        'd1060 :data = 'd1;
        'd1061 :data = 'd0;
        'd1062 :data = 'd1;
        'd1063 :data = 'd0;
        'd1064 :data = 'd0;
        'd1065 :data = 'd0;
        'd1066 :data = 'd1;
        'd1067 :data = 'd1;
        'd1068 :data = 'd1;
        'd1069 :data = 'd1;
        'd1070 :data = 'd0;
        'd1071 :data = 'd0;
        'd1072 :data = 'd1;
        'd1073 :data = 'd1;
        'd1074 :data = 'd1;
        'd1075 :data = 'd0;
        'd1076 :data = 'd0;
        'd1077 :data = 'd1;
        'd1078 :data = 'd0;
        'd1079 :data = 'd0;
        'd1080 :data = 'd0;
        'd1081 :data = 'd1;
        'd1082 :data = 'd0;
        'd1083 :data = 'd1;
        'd1084 :data = 'd1;
        'd1085 :data = 'd0;
        'd1086 :data = 'd0;
        'd1087 :data = 'd0;
        'd1088 :data = 'd0;
        'd1089 :data = 'd0;
        'd1090 :data = 'd0;
        'd1091 :data = 'd1;
        'd1092 :data = 'd1;
        'd1093 :data = 'd1;
        'd1094 :data = 'd1;
        'd1095 :data = 'd0;
        'd1096 :data = 'd0;
        'd1097 :data = 'd1;
        'd1098 :data = 'd1;
        'd1099 :data = 'd1;
        'd1100 :data = 'd0;
        'd1101 :data = 'd1;
        'd1102 :data = 'd1;
        'd1103 :data = 'd1;
        'd1104 :data = 'd0;
        'd1105 :data = 'd0;
        'd1106 :data = 'd0;
        'd1107 :data = 'd1;
        'd1108 :data = 'd1;
        'd1109 :data = 'd1;
        'd1110 :data = 'd0;
        'd1111 :data = 'd1;
        'd1112 :data = 'd0;
        'd1113 :data = 'd0;
        'd1114 :data = 'd0;
        'd1115 :data = 'd0;
        'd1116 :data = 'd1;
        'd1117 :data = 'd0;
        'd1118 :data = 'd0;
        'd1119 :data = 'd0;
        'd1120 :data = 'd1;
        'd1121 :data = 'd0;
        'd1122 :data = 'd1;
        'd1123 :data = 'd0;
        'd1124 :data = 'd1;
        'd1125 :data = 'd0;
        'd1126 :data = 'd1;
        'd1127 :data = 'd1;
        'd1128 :data = 'd1;
        'd1129 :data = 'd1;
        'd1130 :data = 'd1;
        'd1131 :data = 'd0;
        'd1132 :data = 'd1;
        'd1133 :data = 'd1;
        'd1134 :data = 'd0;
        'd1135 :data = 'd1;
        'd1136 :data = 'd0;
        'd1137 :data = 'd0;
        'd1138 :data = 'd0;
        'd1139 :data = 'd1;
        'd1140 :data = 'd1;
        'd1141 :data = 'd1;
        'd1142 :data = 'd0;
        'd1143 :data = 'd1;
        'd1144 :data = 'd1;
        'd1145 :data = 'd1;
        'd1146 :data = 'd0;
        'd1147 :data = 'd1;
        'd1148 :data = 'd0;
        'd1149 :data = 'd0;
        'd1150 :data = 'd0;
        'd1151 :data = 'd0;
        'd1152 :data = 'd0;
        'd1153 :data = 'd0;
        'd1154 :data = 'd0;
        'd1155 :data = 'd0;
        'd1156 :data = 'd0;
        'd1157 :data = 'd0;
        'd1158 :data = 'd1;
        'd1159 :data = 'd1;
        'd1160 :data = 'd1;
        'd1161 :data = 'd0;
        'd1162 :data = 'd0;
        'd1163 :data = 'd1;
        'd1164 :data = 'd1;
        'd1165 :data = 'd0;
        'd1166 :data = 'd0;
        'd1167 :data = 'd0;
        'd1168 :data = 'd1;
        'd1169 :data = 'd1;
        'd1170 :data = 'd1;
        'd1171 :data = 'd1;
        'd1172 :data = 'd1;
        'd1173 :data = 'd0;
        'd1174 :data = 'd1;
        'd1175 :data = 'd0;
        'd1176 :data = 'd1;
        'd1177 :data = 'd0;
        'd1178 :data = 'd1;
        'd1179 :data = 'd1;
        'd1180 :data = 'd1;
        'd1181 :data = 'd0;
        'd1182 :data = 'd0;
        'd1183 :data = 'd0;
        'd1184 :data = 'd0;
        'd1185 :data = 'd0;
        'd1186 :data = 'd0;
        'd1187 :data = 'd0;
        'd1188 :data = 'd0;
        'd1189 :data = 'd0;
        'd1190 :data = 'd1;
        'd1191 :data = 'd1;
        'd1192 :data = 'd1;
        'd1193 :data = 'd0;
        'd1194 :data = 'd0;
        'd1195 :data = 'd0;
        'd1196 :data = 'd0;
        'd1197 :data = 'd1;
        'd1198 :data = 'd1;
        'd1199 :data = 'd0;
        'd1200 :data = 'd0;
        'd1201 :data = 'd0;
        'd1202 :data = 'd0;
        'd1203 :data = 'd0;
        'd1204 :data = 'd1;
        'd1205 :data = 'd0;
        'd1206 :data = 'd0;
        'd1207 :data = 'd1;
        'd1208 :data = 'd0;
        'd1209 :data = 'd0;
        'd1210 :data = 'd0;
        'd1211 :data = 'd1;
        'd1212 :data = 'd1;
        'd1213 :data = 'd0;
        'd1214 :data = 'd0;
        'd1215 :data = 'd1;
        'd1216 :data = 'd0;
        'd1217 :data = 'd1;
        'd1218 :data = 'd1;
        'd1219 :data = 'd1;
        'd1220 :data = 'd1;
        'd1221 :data = 'd0;
        'd1222 :data = 'd1;
        'd1223 :data = 'd0;
        'd1224 :data = 'd1;
        'd1225 :data = 'd0;
        'd1226 :data = 'd0;
        'd1227 :data = 'd1;
        'd1228 :data = 'd0;
        'd1229 :data = 'd0;
        'd1230 :data = 'd1;
        'd1231 :data = 'd0;
        'd1232 :data = 'd1;
        'd1233 :data = 'd0;
        'd1234 :data = 'd1;
        'd1235 :data = 'd0;
        'd1236 :data = 'd0;
        'd1237 :data = 'd0;
        'd1238 :data = 'd1;
        'd1239 :data = 'd1;
        'd1240 :data = 'd1;
        'd1241 :data = 'd0;
        'd1242 :data = 'd0;
        'd1243 :data = 'd0;
        'd1244 :data = 'd1;
        'd1245 :data = 'd0;
        'd1246 :data = 'd1;
        'd1247 :data = 'd0;
        'd1248 :data = 'd0;
        'd1249 :data = 'd1;
        'd1250 :data = 'd1;
        'd1251 :data = 'd1;
        'd1252 :data = 'd0;
        'd1253 :data = 'd1;
        'd1254 :data = 'd1;
        'd1255 :data = 'd0;
        'd1256 :data = 'd0;
        'd1257 :data = 'd1;
        'd1258 :data = 'd1;
        'd1259 :data = 'd0;
        'd1260 :data = 'd0;
        'd1261 :data = 'd0;
        'd1262 :data = 'd0;
        'd1263 :data = 'd0;
        'd1264 :data = 'd1;
        'd1265 :data = 'd0;
        'd1266 :data = 'd1;
        'd1267 :data = 'd1;
        'd1268 :data = 'd0;
        'd1269 :data = 'd0;
        'd1270 :data = 'd0;
        'd1271 :data = 'd0;
        'd1272 :data = 'd1;
        'd1273 :data = 'd1;
        'd1274 :data = 'd0;
        'd1275 :data = 'd1;
        'd1276 :data = 'd1;
        'd1277 :data = 'd1;
        'd1278 :data = 'd0;
        'd1279 :data = 'd0;
        'd1280 :data = 'd0;
        'd1281 :data = 'd1;
        'd1282 :data = 'd0;
        'd1283 :data = 'd0;
        'd1284 :data = 'd1;
        'd1285 :data = 'd1;
        'd1286 :data = 'd1;
        'd1287 :data = 'd1;
        'd1288 :data = 'd1;
        'd1289 :data = 'd0;
        'd1290 :data = 'd0;
        'd1291 :data = 'd0;
        'd1292 :data = 'd0;
        'd1293 :data = 'd0;
        'd1294 :data = 'd1;
        'd1295 :data = 'd0;
        'd1296 :data = 'd0;
        'd1297 :data = 'd0;
        'd1298 :data = 'd0;
        'd1299 :data = 'd0;
        'd1300 :data = 'd0;
        'd1301 :data = 'd1;
        'd1302 :data = 'd0;
        'd1303 :data = 'd0;
        'd1304 :data = 'd1;
        'd1305 :data = 'd0;
        'd1306 :data = 'd1;
        'd1307 :data = 'd0;
        'd1308 :data = 'd1;
        'd1309 :data = 'd0;
        'd1310 :data = 'd0;
        'd1311 :data = 'd0;
        'd1312 :data = 'd1;
        'd1313 :data = 'd0;
        'd1314 :data = 'd0;
        'd1315 :data = 'd0;
        'd1316 :data = 'd0;
        'd1317 :data = 'd0;
        'd1318 :data = 'd0;
        'd1319 :data = 'd1;
        'd1320 :data = 'd1;
        'd1321 :data = 'd1;
        'd1322 :data = 'd1;
        'd1323 :data = 'd0;
        'd1324 :data = 'd1;
        'd1325 :data = 'd0;
        'd1326 :data = 'd1;
        'd1327 :data = 'd1;
        'd1328 :data = 'd0;
        'd1329 :data = 'd0;
        'd1330 :data = 'd1;
        'd1331 :data = 'd0;
        'd1332 :data = 'd0;
        'd1333 :data = 'd0;
        'd1334 :data = 'd0;
        'd1335 :data = 'd1;
        'd1336 :data = 'd1;
        'd1337 :data = 'd0;
        'd1338 :data = 'd1;
        'd1339 :data = 'd1;
        'd1340 :data = 'd1;
        'd1341 :data = 'd0;
        'd1342 :data = 'd1;
        'd1343 :data = 'd0;
        'd1344 :data = 'd1;
        'd1345 :data = 'd0;
        'd1346 :data = 'd0;
        'd1347 :data = 'd0;
        'd1348 :data = 'd1;
        'd1349 :data = 'd1;
        'd1350 :data = 'd0;
        'd1351 :data = 'd1;
        'd1352 :data = 'd1;
        'd1353 :data = 'd0;
        'd1354 :data = 'd0;
        'd1355 :data = 'd0;
        'd1356 :data = 'd1;
        'd1357 :data = 'd0;
        'd1358 :data = 'd1;
        'd1359 :data = 'd0;
        'd1360 :data = 'd0;
        'd1361 :data = 'd0;
        'd1362 :data = 'd0;
        'd1363 :data = 'd1;
        'd1364 :data = 'd1;
        'd1365 :data = 'd1;
        'd1366 :data = 'd0;
        'd1367 :data = 'd1;
        'd1368 :data = 'd0;
        'd1369 :data = 'd0;
        'd1370 :data = 'd1;
        'd1371 :data = 'd1;
        'd1372 :data = 'd0;
        'd1373 :data = 'd0;
        'd1374 :data = 'd1;
        'd1375 :data = 'd0;
        'd1376 :data = 'd0;
        'd1377 :data = 'd0;
        'd1378 :data = 'd0;
        'd1379 :data = 'd1;
        'd1380 :data = 'd1;
        'd1381 :data = 'd0;
        'd1382 :data = 'd1;
        'd1383 :data = 'd1;
        'd1384 :data = 'd1;
        'd1385 :data = 'd1;
        'd1386 :data = 'd0;
        'd1387 :data = 'd0;
        'd1388 :data = 'd0;
        'd1389 :data = 'd1;
        'd1390 :data = 'd1;
        'd1391 :data = 'd1;
        'd1392 :data = 'd1;
        'd1393 :data = 'd1;
        'd1394 :data = 'd1;
        'd1395 :data = 'd1;
        'd1396 :data = 'd0;
        'd1397 :data = 'd0;
        'd1398 :data = 'd0;
        'd1399 :data = 'd1;
        'd1400 :data = 'd0;
        'd1401 :data = 'd1;
        'd1402 :data = 'd1;
        'd1403 :data = 'd0;
        'd1404 :data = 'd0;
        'd1405 :data = 'd1;
        'd1406 :data = 'd1;
        'd1407 :data = 'd1;
        'd1408 :data = 'd0;
        'd1409 :data = 'd1;
        'd1410 :data = 'd1;
        'd1411 :data = 'd1;
        'd1412 :data = 'd1;
        'd1413 :data = 'd1;
        'd1414 :data = 'd0;
        'd1415 :data = 'd1;
        'd1416 :data = 'd1;
        'd1417 :data = 'd1;
        'd1418 :data = 'd1;
        'd1419 :data = 'd0;
        'd1420 :data = 'd1;
        'd1421 :data = 'd1;
        'd1422 :data = 'd0;
        'd1423 :data = 'd0;
        'd1424 :data = 'd0;
        'd1425 :data = 'd0;
        'd1426 :data = 'd0;
        'd1427 :data = 'd0;
        'd1428 :data = 'd0;
        'd1429 :data = 'd0;
        'd1430 :data = 'd0;
        'd1431 :data = 'd0;
        'd1432 :data = 'd1;
        'd1433 :data = 'd0;
        'd1434 :data = 'd0;
        'd1435 :data = 'd1;
        'd1436 :data = 'd1;
        'd1437 :data = 'd0;
        'd1438 :data = 'd0;
        'd1439 :data = 'd0;
        'd1440 :data = 'd1;
        'd1441 :data = 'd1;
        'd1442 :data = 'd1;
        'd1443 :data = 'd0;
        'd1444 :data = 'd0;
        'd1445 :data = 'd1;
        'd1446 :data = 'd1;
        'd1447 :data = 'd0;
        'd1448 :data = 'd0;
        'd1449 :data = 'd1;
        'd1450 :data = 'd0;
        'd1451 :data = 'd0;
        'd1452 :data = 'd1;
        'd1453 :data = 'd0;
        'd1454 :data = 'd1;
        'd1455 :data = 'd1;
        'd1456 :data = 'd1;
        'd1457 :data = 'd0;
        'd1458 :data = 'd0;
        'd1459 :data = 'd1;
        'd1460 :data = 'd0;
        'd1461 :data = 'd1;
        'd1462 :data = 'd0;
        'd1463 :data = 'd1;
        'd1464 :data = 'd0;
        'd1465 :data = 'd0;
        'd1466 :data = 'd1;
        'd1467 :data = 'd1;
        'd1468 :data = 'd0;
        'd1469 :data = 'd0;
        'd1470 :data = 'd0;
        'd1471 :data = 'd1;
        'd1472 :data = 'd0;
        'd1473 :data = 'd0;
        'd1474 :data = 'd0;
        'd1475 :data = 'd0;
        'd1476 :data = 'd1;
        'd1477 :data = 'd0;
        'd1478 :data = 'd0;
        'd1479 :data = 'd0;
        'd1480 :data = 'd0;
        'd1481 :data = 'd0;
        'd1482 :data = 'd0;
        'd1483 :data = 'd0;
        'd1484 :data = 'd1;
        'd1485 :data = 'd1;
        'd1486 :data = 'd1;
        'd1487 :data = 'd0;
        'd1488 :data = 'd1;
        'd1489 :data = 'd0;
        'd1490 :data = 'd1;
        'd1491 :data = 'd0;
        'd1492 :data = 'd0;
        'd1493 :data = 'd0;
        'd1494 :data = 'd0;
        'd1495 :data = 'd0;
        'd1496 :data = 'd1;
        'd1497 :data = 'd0;
        'd1498 :data = 'd0;
        'd1499 :data = 'd0;
        'd1500 :data = 'd1;
        'd1501 :data = 'd1;
        'd1502 :data = 'd1;
        'd1503 :data = 'd1;
        'd1504 :data = 'd0;
        'd1505 :data = 'd0;
        'd1506 :data = 'd1;
        'd1507 :data = 'd1;
        'd1508 :data = 'd0;
        'd1509 :data = 'd0;
        'd1510 :data = 'd0;
        'd1511 :data = 'd0;
        'd1512 :data = 'd0;
        'd1513 :data = 'd0;
        'd1514 :data = 'd0;
        'd1515 :data = 'd1;
        'd1516 :data = 'd0;
        'd1517 :data = 'd0;
        'd1518 :data = 'd0;
        'd1519 :data = 'd1;
        'd1520 :data = 'd0;
        'd1521 :data = 'd1;
        'd1522 :data = 'd1;
        'd1523 :data = 'd1;
        'd1524 :data = 'd1;
        'd1525 :data = 'd1;
        'd1526 :data = 'd0;
        'd1527 :data = 'd1;
        'd1528 :data = 'd1;
        'd1529 :data = 'd0;
        'd1530 :data = 'd0;
        'd1531 :data = 'd0;
        'd1532 :data = 'd0;
        'd1533 :data = 'd0;
        'd1534 :data = 'd0;
        'd1535 :data = 'd0;
        'd1536 :data = 'd0;
        'd1537 :data = 'd0;
        'd1538 :data = 'd1;
        'd1539 :data = 'd0;
        'd1540 :data = 'd0;
        'd1541 :data = 'd0;
        'd1542 :data = 'd0;
        'd1543 :data = 'd0;
        'd1544 :data = 'd0;
        'd1545 :data = 'd1;
        'd1546 :data = 'd1;
        'd1547 :data = 'd0;
        'd1548 :data = 'd0;
        'd1549 :data = 'd0;
        'd1550 :data = 'd1;
        'd1551 :data = 'd1;
        'd1552 :data = 'd0;
        'd1553 :data = 'd0;
        'd1554 :data = 'd0;
        'd1555 :data = 'd1;
        'd1556 :data = 'd1;
        'd1557 :data = 'd1;
        'd1558 :data = 'd0;
        'd1559 :data = 'd1;
        'd1560 :data = 'd1;
        'd1561 :data = 'd0;
        'd1562 :data = 'd1;
        'd1563 :data = 'd1;
        'd1564 :data = 'd0;
        'd1565 :data = 'd0;
        'd1566 :data = 'd1;
        'd1567 :data = 'd1;
        'd1568 :data = 'd1;
        'd1569 :data = 'd0;
        'd1570 :data = 'd0;
        'd1571 :data = 'd1;
        'd1572 :data = 'd1;
        'd1573 :data = 'd0;
        'd1574 :data = 'd0;
        'd1575 :data = 'd0;
        'd1576 :data = 'd1;
        'd1577 :data = 'd1;
        'd1578 :data = 'd1;
        'd1579 :data = 'd1;
        'd1580 :data = 'd0;
        'd1581 :data = 'd0;
        'd1582 :data = 'd0;
        'd1583 :data = 'd0;
        'd1584 :data = 'd1;
        'd1585 :data = 'd1;
        'd1586 :data = 'd1;
        'd1587 :data = 'd0;
        'd1588 :data = 'd0;
        'd1589 :data = 'd1;
        'd1590 :data = 'd0;
        'd1591 :data = 'd0;
        'd1592 :data = 'd0;
        'd1593 :data = 'd1;
        'd1594 :data = 'd1;
        'd1595 :data = 'd0;
        'd1596 :data = 'd0;
        'd1597 :data = 'd1;
        'd1598 :data = 'd0;
        'd1599 :data = 'd1;
        'd1600 :data = 'd1;
        'd1601 :data = 'd0;
        'd1602 :data = 'd1;
        'd1603 :data = 'd0;
        'd1604 :data = 'd0;
        'd1605 :data = 'd1;
        'd1606 :data = 'd1;
        'd1607 :data = 'd0;
        'd1608 :data = 'd0;
        'd1609 :data = 'd1;
        'd1610 :data = 'd1;
        'd1611 :data = 'd0;
        'd1612 :data = 'd1;
        'd1613 :data = 'd1;
        'd1614 :data = 'd0;
        'd1615 :data = 'd0;
        'd1616 :data = 'd1;
        'd1617 :data = 'd0;
        'd1618 :data = 'd1;
        'd1619 :data = 'd1;
        'd1620 :data = 'd1;
        'd1621 :data = 'd1;
        'd1622 :data = 'd0;
        'd1623 :data = 'd1;
        'd1624 :data = 'd0;
        'd1625 :data = 'd1;
        'd1626 :data = 'd1;
        'd1627 :data = 'd1;
        'd1628 :data = 'd1;
        'd1629 :data = 'd1;
        'd1630 :data = 'd1;
        'd1631 :data = 'd1;
        'd1632 :data = 'd0;
        'd1633 :data = 'd1;
        'd1634 :data = 'd1;
        'd1635 :data = 'd1;
        'd1636 :data = 'd0;
        'd1637 :data = 'd0;
        'd1638 :data = 'd0;
        'd1639 :data = 'd0;
        'd1640 :data = 'd0;
        'd1641 :data = 'd1;
        'd1642 :data = 'd0;
        'd1643 :data = 'd0;
        'd1644 :data = 'd1;
        'd1645 :data = 'd0;
        'd1646 :data = 'd1;
        'd1647 :data = 'd0;
        'd1648 :data = 'd0;
        'd1649 :data = 'd0;
        'd1650 :data = 'd1;
        'd1651 :data = 'd0;
        'd1652 :data = 'd0;
        'd1653 :data = 'd0;
        'd1654 :data = 'd0;
        'd1655 :data = 'd0;
        'd1656 :data = 'd0;
        'd1657 :data = 'd1;
        'd1658 :data = 'd0;
        'd1659 :data = 'd1;
        'd1660 :data = 'd1;
        'd1661 :data = 'd1;
        'd1662 :data = 'd1;
        'd1663 :data = 'd0;
        'd1664 :data = 'd0;
        'd1665 :data = 'd0;
        'd1666 :data = 'd0;
        'd1667 :data = 'd1;
        'd1668 :data = 'd1;
        'd1669 :data = 'd1;
        'd1670 :data = 'd0;
        'd1671 :data = 'd1;
        'd1672 :data = 'd0;
        'd1673 :data = 'd1;
        'd1674 :data = 'd0;
        'd1675 :data = 'd0;
        'd1676 :data = 'd1;
        'd1677 :data = 'd0;
        'd1678 :data = 'd1;
        'd1679 :data = 'd1;
        'd1680 :data = 'd0;
        'd1681 :data = 'd1;
        'd1682 :data = 'd0;
        'd1683 :data = 'd0;
        'd1684 :data = 'd1;
        'd1685 :data = 'd1;
        'd1686 :data = 'd1;
        'd1687 :data = 'd0;
        'd1688 :data = 'd1;
        'd1689 :data = 'd0;
        'd1690 :data = 'd1;
        'd1691 :data = 'd0;
        'd1692 :data = 'd1;
        'd1693 :data = 'd0;
        'd1694 :data = 'd1;
        'd1695 :data = 'd0;
        'd1696 :data = 'd1;
        'd1697 :data = 'd0;
        'd1698 :data = 'd0;
        'd1699 :data = 'd0;
        'd1700 :data = 'd0;
        'd1701 :data = 'd0;
        'd1702 :data = 'd1;
        'd1703 :data = 'd1;
        'd1704 :data = 'd0;
        'd1705 :data = 'd0;
        'd1706 :data = 'd0;
        'd1707 :data = 'd1;
        'd1708 :data = 'd1;
        'd1709 :data = 'd1;
        'd1710 :data = 'd0;
        'd1711 :data = 'd1;
        'd1712 :data = 'd0;
        'd1713 :data = 'd1;
        'd1714 :data = 'd1;
        'd1715 :data = 'd0;
        'd1716 :data = 'd0;
        'd1717 :data = 'd0;
        'd1718 :data = 'd1;
        'd1719 :data = 'd0;
        'd1720 :data = 'd0;
        'd1721 :data = 'd1;
        'd1722 :data = 'd0;
        'd1723 :data = 'd0;
        'd1724 :data = 'd0;
        'd1725 :data = 'd0;
        'd1726 :data = 'd1;
        'd1727 :data = 'd1;
        'd1728 :data = 'd0;
        'd1729 :data = 'd0;
        'd1730 :data = 'd0;
        'd1731 :data = 'd0;
        'd1732 :data = 'd0;
        'd1733 :data = 'd1;
        'd1734 :data = 'd1;
        'd1735 :data = 'd0;
        'd1736 :data = 'd1;
        'd1737 :data = 'd0;
        'd1738 :data = 'd1;
        'd1739 :data = 'd1;
        'd1740 :data = 'd0;
        'd1741 :data = 'd1;
        'd1742 :data = 'd1;
        'd1743 :data = 'd0;
        'd1744 :data = 'd1;
        'd1745 :data = 'd0;
        'd1746 :data = 'd0;
        'd1747 :data = 'd1;
        'd1748 :data = 'd1;
        'd1749 :data = 'd1;
        'd1750 :data = 'd1;
        'd1751 :data = 'd0;
        'd1752 :data = 'd1;
        'd1753 :data = 'd1;
        'd1754 :data = 'd1;
        'd1755 :data = 'd0;
        'd1756 :data = 'd0;
        'd1757 :data = 'd0;
        'd1758 :data = 'd1;
        'd1759 :data = 'd0;
        'd1760 :data = 'd0;
        'd1761 :data = 'd0;
        'd1762 :data = 'd0;
        'd1763 :data = 'd1;
        'd1764 :data = 'd1;
        'd1765 :data = 'd0;
        'd1766 :data = 'd0;
        'd1767 :data = 'd0;
        'd1768 :data = 'd1;
        'd1769 :data = 'd1;
        'd1770 :data = 'd1;
        'd1771 :data = 'd1;
        'd1772 :data = 'd1;
        'd1773 :data = 'd1;
        'd1774 :data = 'd1;
        'd1775 :data = 'd1;
        'd1776 :data = 'd1;
        'd1777 :data = 'd0;
        'd1778 :data = 'd0;
        'd1779 :data = 'd1;
        'd1780 :data = 'd1;
        'd1781 :data = 'd1;
        'd1782 :data = 'd1;
        'd1783 :data = 'd0;
        'd1784 :data = 'd1;
        'd1785 :data = 'd1;
        'd1786 :data = 'd1;
        'd1787 :data = 'd0;
        'd1788 :data = 'd0;
        'd1789 :data = 'd1;
        'd1790 :data = 'd1;
        'd1791 :data = 'd0;
        'd1792 :data = 'd1;
        'd1793 :data = 'd1;
        'd1794 :data = 'd1;
        'd1795 :data = 'd0;
        'd1796 :data = 'd0;
        'd1797 :data = 'd0;
        'd1798 :data = 'd0;
        'd1799 :data = 'd0;
        'd1800 :data = 'd0;
        'd1801 :data = 'd0;
        'd1802 :data = 'd1;
        'd1803 :data = 'd0;
        'd1804 :data = 'd1;
        'd1805 :data = 'd1;
        'd1806 :data = 'd1;
        'd1807 :data = 'd1;
        'd1808 :data = 'd0;
        'd1809 :data = 'd0;
        'd1810 :data = 'd0;
        'd1811 :data = 'd1;
        'd1812 :data = 'd1;
        'd1813 :data = 'd1;
        'd1814 :data = 'd1;
        'd1815 :data = 'd1;
        'd1816 :data = 'd1;
        'd1817 :data = 'd1;
        'd1818 :data = 'd0;
        'd1819 :data = 'd1;
        'd1820 :data = 'd0;
        'd1821 :data = 'd1;
        'd1822 :data = 'd0;
        'd1823 :data = 'd1;
        'd1824 :data = 'd0;
        'd1825 :data = 'd0;
        'd1826 :data = 'd1;
        'd1827 :data = 'd0;
        'd1828 :data = 'd0;
        'd1829 :data = 'd0;
        'd1830 :data = 'd0;
        'd1831 :data = 'd0;
        'd1832 :data = 'd0;
        'd1833 :data = 'd0;
        'd1834 :data = 'd0;
        'd1835 :data = 'd1;
        'd1836 :data = 'd1;
        'd1837 :data = 'd1;
        'd1838 :data = 'd0;
        'd1839 :data = 'd0;
        'd1840 :data = 'd0;
        'd1841 :data = 'd0;
        'd1842 :data = 'd0;
        'd1843 :data = 'd1;
        'd1844 :data = 'd0;
        'd1845 :data = 'd1;
        'd1846 :data = 'd1;
        'd1847 :data = 'd1;
        'd1848 :data = 'd1;
        'd1849 :data = 'd1;
        'd1850 :data = 'd0;
        'd1851 :data = 'd1;
        'd1852 :data = 'd0;
        'd1853 :data = 'd0;
        'd1854 :data = 'd1;
        'd1855 :data = 'd0;
        'd1856 :data = 'd0;
        'd1857 :data = 'd0;
        'd1858 :data = 'd0;
        'd1859 :data = 'd0;
        'd1860 :data = 'd1;
        'd1861 :data = 'd1;
        'd1862 :data = 'd1;
        'd1863 :data = 'd0;
        'd1864 :data = 'd1;
        'd1865 :data = 'd0;
        'd1866 :data = 'd1;
        'd1867 :data = 'd0;
        'd1868 :data = 'd1;
        'd1869 :data = 'd0;
        'd1870 :data = 'd1;
        'd1871 :data = 'd1;
        'd1872 :data = 'd1;
        'd1873 :data = 'd0;
        'd1874 :data = 'd1;
        'd1875 :data = 'd0;
        'd1876 :data = 'd1;
        'd1877 :data = 'd1;
        'd1878 :data = 'd1;
        'd1879 :data = 'd1;
        'd1880 :data = 'd1;
        'd1881 :data = 'd0;
        'd1882 :data = 'd0;
        'd1883 :data = 'd1;
        'd1884 :data = 'd0;
        'd1885 :data = 'd1;
        'd1886 :data = 'd0;
        'd1887 :data = 'd0;
        'd1888 :data = 'd0;
        'd1889 :data = 'd0;
        'd1890 :data = 'd0;
        'd1891 :data = 'd1;
        'd1892 :data = 'd0;
        'd1893 :data = 'd1;
        'd1894 :data = 'd0;
        'd1895 :data = 'd0;
        'd1896 :data = 'd1;
        'd1897 :data = 'd1;
        'd1898 :data = 'd0;
        'd1899 :data = 'd0;
        'd1900 :data = 'd0;
        'd1901 :data = 'd1;
        'd1902 :data = 'd1;
        'd1903 :data = 'd1;
        'd1904 :data = 'd0;
        'd1905 :data = 'd1;
        'd1906 :data = 'd0;
        'd1907 :data = 'd1;
        'd1908 :data = 'd0;
        'd1909 :data = 'd1;
        'd1910 :data = 'd0;
        'd1911 :data = 'd0;
        'd1912 :data = 'd1;
        'd1913 :data = 'd1;
        'd1914 :data = 'd0;
        'd1915 :data = 'd1;
        'd1916 :data = 'd0;
        'd1917 :data = 'd1;
        'd1918 :data = 'd1;
        'd1919 :data = 'd1;
        'd1920 :data = 'd0;
        'd1921 :data = 'd1;
        'd1922 :data = 'd0;
        'd1923 :data = 'd0;
        'd1924 :data = 'd1;
        'd1925 :data = 'd1;
        'd1926 :data = 'd0;
        'd1927 :data = 'd1;
        'd1928 :data = 'd0;
        'd1929 :data = 'd1;
        'd1930 :data = 'd1;
        'd1931 :data = 'd1;
        'd1932 :data = 'd1;
        'd1933 :data = 'd0;
        'd1934 :data = 'd1;
        'd1935 :data = 'd0;
        'd1936 :data = 'd1;
        'd1937 :data = 'd1;
        'd1938 :data = 'd0;
        'd1939 :data = 'd1;
        'd1940 :data = 'd0;
        'd1941 :data = 'd1;
        'd1942 :data = 'd1;
        'd1943 :data = 'd0;
        'd1944 :data = 'd1;
        'd1945 :data = 'd1;
        'd1946 :data = 'd0;
        'd1947 :data = 'd0;
        'd1948 :data = 'd0;
        'd1949 :data = 'd0;
        'd1950 :data = 'd1;
        'd1951 :data = 'd0;
        'd1952 :data = 'd0;
        'd1953 :data = 'd1;
        'd1954 :data = 'd0;
        'd1955 :data = 'd0;
        'd1956 :data = 'd1;
        'd1957 :data = 'd1;
        'd1958 :data = 'd1;
        'd1959 :data = 'd0;
        'd1960 :data = 'd0;
        'd1961 :data = 'd1;
        'd1962 :data = 'd0;
        'd1963 :data = 'd1;
        'd1964 :data = 'd1;
        'd1965 :data = 'd1;
        'd1966 :data = 'd1;
        'd1967 :data = 'd0;
        'd1968 :data = 'd1;
        'd1969 :data = 'd0;
        'd1970 :data = 'd0;
        'd1971 :data = 'd1;
        'd1972 :data = 'd1;
        'd1973 :data = 'd1;
        'd1974 :data = 'd1;
        'd1975 :data = 'd0;
        'd1976 :data = 'd1;
        'd1977 :data = 'd1;
        'd1978 :data = 'd1;
        'd1979 :data = 'd1;
        'd1980 :data = 'd0;
        'd1981 :data = 'd0;
        'd1982 :data = 'd0;
        'd1983 :data = 'd0;
        'd1984 :data = 'd0;
        'd1985 :data = 'd0;
        'd1986 :data = 'd1;
        'd1987 :data = 'd1;
        'd1988 :data = 'd1;
        'd1989 :data = 'd0;
        'd1990 :data = 'd1;
        'd1991 :data = 'd0;
        'd1992 :data = 'd0;
        'd1993 :data = 'd0;
        'd1994 :data = 'd1;
        'd1995 :data = 'd0;
        'd1996 :data = 'd1;
        'd1997 :data = 'd1;
        'd1998 :data = 'd1;
        'd1999 :data = 'd1;
        'd2000 :data = 'd0;
        'd2001 :data = 'd0;
        'd2002 :data = 'd1;
        'd2003 :data = 'd1;
        'd2004 :data = 'd0;
        'd2005 :data = 'd0;
        'd2006 :data = 'd1;
        'd2007 :data = 'd0;
        'd2008 :data = 'd1;
        'd2009 :data = 'd0;
        'd2010 :data = 'd1;
        'd2011 :data = 'd0;
        'd2012 :data = 'd1;
        'd2013 :data = 'd1;
        'd2014 :data = 'd0;
        'd2015 :data = 'd1;
        'd2016 :data = 'd1;
        'd2017 :data = 'd0;
        'd2018 :data = 'd0;
        'd2019 :data = 'd1;
        'd2020 :data = 'd0;
        'd2021 :data = 'd1;
        'd2022 :data = 'd1;
        'd2023 :data = 'd1;
        'd2024 :data = 'd1;
        'd2025 :data = 'd0;
        'd2026 :data = 'd1;
        'd2027 :data = 'd1;
        'd2028 :data = 'd1;
        'd2029 :data = 'd0;
        'd2030 :data = 'd0;
        'd2031 :data = 'd0;
        'd2032 :data = 'd0;
        'd2033 :data = 'd1;
        'd2034 :data = 'd1;
        'd2035 :data = 'd1;
        'd2036 :data = 'd1;
        'd2037 :data = 'd1;
        'd2038 :data = 'd0;
        'd2039 :data = 'd1;
        'd2040 :data = 'd0;
        'd2041 :data = 'd0;
        'd2042 :data = 'd0;
        'd2043 :data = 'd0;
        'd2044 :data = 'd1;
        'd2045 :data = 'd1;
        'd2046 :data = 'd1;
        'd2047 :data = 'd0;
        'd2048 :data = 'd0;
        'd2049 :data = 'd0;
        'd2050 :data = 'd1;
        'd2051 :data = 'd1;
        'd2052 :data = 'd1;
        'd2053 :data = 'd1;
        'd2054 :data = 'd1;
        'd2055 :data = 'd1;
        'd2056 :data = 'd1;
        'd2057 :data = 'd0;
        'd2058 :data = 'd1;
        'd2059 :data = 'd0;
        'd2060 :data = 'd0;
        'd2061 :data = 'd0;
        'd2062 :data = 'd1;
        'd2063 :data = 'd1;
        'd2064 :data = 'd0;
        'd2065 :data = 'd0;
        'd2066 :data = 'd0;
        'd2067 :data = 'd0;
        'd2068 :data = 'd0;
        'd2069 :data = 'd1;
        'd2070 :data = 'd0;
        'd2071 :data = 'd0;
        'd2072 :data = 'd0;
        'd2073 :data = 'd1;
        'd2074 :data = 'd1;
        'd2075 :data = 'd1;
        'd2076 :data = 'd0;
        'd2077 :data = 'd1;
        'd2078 :data = 'd1;
        'd2079 :data = 'd0;
        'd2080 :data = 'd1;
        'd2081 :data = 'd1;
        'd2082 :data = 'd0;
        'd2083 :data = 'd1;
        'd2084 :data = 'd0;
        'd2085 :data = 'd0;
        'd2086 :data = 'd0;
        'd2087 :data = 'd1;
        'd2088 :data = 'd1;
        'd2089 :data = 'd1;
        'd2090 :data = 'd0;
        'd2091 :data = 'd0;
        'd2092 :data = 'd0;
        'd2093 :data = 'd1;
        'd2094 :data = 'd0;
        'd2095 :data = 'd1;
        'd2096 :data = 'd0;
        'd2097 :data = 'd0;
        'd2098 :data = 'd0;
        'd2099 :data = 'd1;
        'd2100 :data = 'd0;
        'd2101 :data = 'd0;
        'd2102 :data = 'd0;
        'd2103 :data = 'd1;
        'd2104 :data = 'd1;
        'd2105 :data = 'd1;
        'd2106 :data = 'd1;
        'd2107 :data = 'd1;
        'd2108 :data = 'd0;
        'd2109 :data = 'd0;
        'd2110 :data = 'd1;
        'd2111 :data = 'd0;
        'd2112 :data = 'd1;
        'd2113 :data = 'd0;
        'd2114 :data = 'd1;
        'd2115 :data = 'd0;
        'd2116 :data = 'd1;
        'd2117 :data = 'd0;
        'd2118 :data = 'd0;
        'd2119 :data = 'd1;
        'd2120 :data = 'd1;
        'd2121 :data = 'd1;
        'd2122 :data = 'd0;
        'd2123 :data = 'd1;
        'd2124 :data = 'd0;
        'd2125 :data = 'd0;
        'd2126 :data = 'd0;
        'd2127 :data = 'd1;
        'd2128 :data = 'd1;
        'd2129 :data = 'd0;
        'd2130 :data = 'd1;
        'd2131 :data = 'd1;
        'd2132 :data = 'd0;
        'd2133 :data = 'd0;
        'd2134 :data = 'd0;
        'd2135 :data = 'd0;
        'd2136 :data = 'd1;
        'd2137 :data = 'd0;
        'd2138 :data = 'd0;
        'd2139 :data = 'd1;
        'd2140 :data = 'd1;
        'd2141 :data = 'd0;
        'd2142 :data = 'd0;
        'd2143 :data = 'd0;
        'd2144 :data = 'd0;
        'd2145 :data = 'd1;
        'd2146 :data = 'd1;
        'd2147 :data = 'd1;
        'd2148 :data = 'd0;
        'd2149 :data = 'd1;
        'd2150 :data = 'd0;
        'd2151 :data = 'd0;
        'd2152 :data = 'd1;
        'd2153 :data = 'd0;
        'd2154 :data = 'd1;
        'd2155 :data = 'd1;
        'd2156 :data = 'd1;
        'd2157 :data = 'd0;
        'd2158 :data = 'd0;
        'd2159 :data = 'd0;
        'd2160 :data = 'd1;
        'd2161 :data = 'd1;
        'd2162 :data = 'd0;
        'd2163 :data = 'd1;
        'd2164 :data = 'd0;
        'd2165 :data = 'd1;
        'd2166 :data = 'd1;
        'd2167 :data = 'd1;
        'd2168 :data = 'd1;
        'd2169 :data = 'd0;
        'd2170 :data = 'd1;
        'd2171 :data = 'd1;
        'd2172 :data = 'd0;
        'd2173 :data = 'd1;
        'd2174 :data = 'd1;
        'd2175 :data = 'd0;
        'd2176 :data = 'd0;
        'd2177 :data = 'd1;
        'd2178 :data = 'd0;
        'd2179 :data = 'd0;
        'd2180 :data = 'd0;
        'd2181 :data = 'd0;
        'd2182 :data = 'd1;
        'd2183 :data = 'd0;
        'd2184 :data = 'd0;
        'd2185 :data = 'd0;
        'd2186 :data = 'd1;
        'd2187 :data = 'd1;
        'd2188 :data = 'd1;
        'd2189 :data = 'd1;
        'd2190 :data = 'd0;
        'd2191 :data = 'd1;
        'd2192 :data = 'd0;
        'd2193 :data = 'd1;
        'd2194 :data = 'd1;
        'd2195 :data = 'd1;
        'd2196 :data = 'd1;
        'd2197 :data = 'd1;
        'd2198 :data = 'd0;
        'd2199 :data = 'd0;
        'd2200 :data = 'd1;
        'd2201 :data = 'd1;
        'd2202 :data = 'd0;
        'd2203 :data = 'd0;
        'd2204 :data = 'd0;
        'd2205 :data = 'd1;
        'd2206 :data = 'd1;
        'd2207 :data = 'd0;
        'd2208 :data = 'd1;
        'd2209 :data = 'd0;
        'd2210 :data = 'd0;
        'd2211 :data = 'd1;
        'd2212 :data = 'd1;
        'd2213 :data = 'd0;
        'd2214 :data = 'd0;
        'd2215 :data = 'd0;
        'd2216 :data = 'd1;
        'd2217 :data = 'd1;
        'd2218 :data = 'd1;
        'd2219 :data = 'd1;
        'd2220 :data = 'd0;
        'd2221 :data = 'd0;
        'd2222 :data = 'd1;
        'd2223 :data = 'd1;
        'd2224 :data = 'd1;
        'd2225 :data = 'd0;
        'd2226 :data = 'd0;
        'd2227 :data = 'd1;
        'd2228 :data = 'd0;
        'd2229 :data = 'd1;
        'd2230 :data = 'd1;
        'd2231 :data = 'd0;
        'd2232 :data = 'd1;
        'd2233 :data = 'd1;
        'd2234 :data = 'd1;
        'd2235 :data = 'd0;
        'd2236 :data = 'd0;
        'd2237 :data = 'd0;
        'd2238 :data = 'd0;
        'd2239 :data = 'd0;
        'd2240 :data = 'd0;
        'd2241 :data = 'd0;
        'd2242 :data = 'd1;
        'd2243 :data = 'd0;
        'd2244 :data = 'd1;
        'd2245 :data = 'd0;
        'd2246 :data = 'd1;
        'd2247 :data = 'd1;
        'd2248 :data = 'd0;
        'd2249 :data = 'd1;
        'd2250 :data = 'd0;
        'd2251 :data = 'd0;
        'd2252 :data = 'd0;
        'd2253 :data = 'd1;
        'd2254 :data = 'd1;
        'd2255 :data = 'd1;
        'd2256 :data = 'd0;
        'd2257 :data = 'd0;
        'd2258 :data = 'd1;
        'd2259 :data = 'd1;
        'd2260 :data = 'd0;
        'd2261 :data = 'd1;
        'd2262 :data = 'd1;
        'd2263 :data = 'd1;
        'd2264 :data = 'd1;
        'd2265 :data = 'd0;
        'd2266 :data = 'd1;
        'd2267 :data = 'd1;
        'd2268 :data = 'd1;
        'd2269 :data = 'd1;
        'd2270 :data = 'd0;
        'd2271 :data = 'd1;
        'd2272 :data = 'd0;
        'd2273 :data = 'd1;
        'd2274 :data = 'd1;
        'd2275 :data = 'd1;
        'd2276 :data = 'd0;
        'd2277 :data = 'd1;
        'd2278 :data = 'd0;
        'd2279 :data = 'd1;
        'd2280 :data = 'd0;
        'd2281 :data = 'd1;
        'd2282 :data = 'd0;
        'd2283 :data = 'd1;
        'd2284 :data = 'd0;
        'd2285 :data = 'd0;
        'd2286 :data = 'd0;
        'd2287 :data = 'd1;
        'd2288 :data = 'd0;
        'd2289 :data = 'd0;
        'd2290 :data = 'd1;
        'd2291 :data = 'd0;
        'd2292 :data = 'd1;
        'd2293 :data = 'd0;
        'd2294 :data = 'd1;
        'd2295 :data = 'd0;
        'd2296 :data = 'd1;
        'd2297 :data = 'd0;
        'd2298 :data = 'd0;
        'd2299 :data = 'd0;
        'd2300 :data = 'd1;
        'd2301 :data = 'd1;
        'd2302 :data = 'd0;
        'd2303 :data = 'd0;
        'd2304 :data = 'd0;
        'd2305 :data = 'd1;
        'd2306 :data = 'd0;
        'd2307 :data = 'd0;
        'd2308 :data = 'd1;
        'd2309 :data = 'd1;
        'd2310 :data = 'd1;
        'd2311 :data = 'd0;
        'd2312 :data = 'd0;
        'd2313 :data = 'd0;
        'd2314 :data = 'd1;
        'd2315 :data = 'd1;
        'd2316 :data = 'd1;
        'd2317 :data = 'd0;
        'd2318 :data = 'd0;
        'd2319 :data = 'd1;
        'd2320 :data = 'd0;
        'd2321 :data = 'd1;
        'd2322 :data = 'd0;
        'd2323 :data = 'd0;
        'd2324 :data = 'd0;
        'd2325 :data = 'd0;
        'd2326 :data = 'd1;
        'd2327 :data = 'd0;
        'd2328 :data = 'd1;
        'd2329 :data = 'd0;
        'd2330 :data = 'd0;
        'd2331 :data = 'd0;
        'd2332 :data = 'd0;
        'd2333 :data = 'd0;
        'd2334 :data = 'd1;
        'd2335 :data = 'd1;
        'd2336 :data = 'd0;
        'd2337 :data = 'd0;
        'd2338 :data = 'd1;
        'd2339 :data = 'd1;
        'd2340 :data = 'd0;
        'd2341 :data = 'd1;
        'd2342 :data = 'd1;
        'd2343 :data = 'd1;
        'd2344 :data = 'd1;
        'd2345 :data = 'd0;
        'd2346 :data = 'd0;
        'd2347 :data = 'd0;
        'd2348 :data = 'd1;
        'd2349 :data = 'd1;
        'd2350 :data = 'd0;
        'd2351 :data = 'd0;
        'd2352 :data = 'd1;
        'd2353 :data = 'd0;
        'd2354 :data = 'd1;
        'd2355 :data = 'd1;
        'd2356 :data = 'd0;
        'd2357 :data = 'd1;
        'd2358 :data = 'd1;
        'd2359 :data = 'd1;
        'd2360 :data = 'd1;
        'd2361 :data = 'd0;
        'd2362 :data = 'd1;
        'd2363 :data = 'd0;
        'd2364 :data = 'd1;
        'd2365 :data = 'd0;
        'd2366 :data = 'd0;
        'd2367 :data = 'd0;
        'd2368 :data = 'd1;
        'd2369 :data = 'd1;
        'd2370 :data = 'd1;
        'd2371 :data = 'd0;
        'd2372 :data = 'd0;
        'd2373 :data = 'd1;
        'd2374 :data = 'd1;
        'd2375 :data = 'd0;
        'd2376 :data = 'd0;
        'd2377 :data = 'd1;
        'd2378 :data = 'd1;
        'd2379 :data = 'd0;
        'd2380 :data = 'd1;
        'd2381 :data = 'd1;
        'd2382 :data = 'd0;
        'd2383 :data = 'd0;
        'd2384 :data = 'd0;
        'd2385 :data = 'd1;
        'd2386 :data = 'd0;
        'd2387 :data = 'd1;
        'd2388 :data = 'd1;
        'd2389 :data = 'd1;
        'd2390 :data = 'd1;
        'd2391 :data = 'd0;
        'd2392 :data = 'd1;
        'd2393 :data = 'd0;
        'd2394 :data = 'd1;
        'd2395 :data = 'd0;
        'd2396 :data = 'd1;
        'd2397 :data = 'd1;
        'd2398 :data = 'd0;
        'd2399 :data = 'd0;
        'd2400 :data = 'd1;
        'd2401 :data = 'd0;
        'd2402 :data = 'd1;
        'd2403 :data = 'd1;
        'd2404 :data = 'd0;
        'd2405 :data = 'd0;
        'd2406 :data = 'd0;
        'd2407 :data = 'd1;
        'd2408 :data = 'd0;
        'd2409 :data = 'd1;
        'd2410 :data = 'd0;
        'd2411 :data = 'd1;
        'd2412 :data = 'd1;
        'd2413 :data = 'd1;
        'd2414 :data = 'd1;
        'd2415 :data = 'd1;
        'd2416 :data = 'd0;
        'd2417 :data = 'd0;
        'd2418 :data = 'd0;
        'd2419 :data = 'd1;
        'd2420 :data = 'd1;
        'd2421 :data = 'd0;
        'd2422 :data = 'd0;
        'd2423 :data = 'd1;
        'd2424 :data = 'd1;
        'd2425 :data = 'd1;
        'd2426 :data = 'd0;
        'd2427 :data = 'd0;
        'd2428 :data = 'd0;
        'd2429 :data = 'd1;
        'd2430 :data = 'd0;
        'd2431 :data = 'd1;
        'd2432 :data = 'd0;
        'd2433 :data = 'd0;
        'd2434 :data = 'd0;
        'd2435 :data = 'd0;
        'd2436 :data = 'd1;
        'd2437 :data = 'd0;
        'd2438 :data = 'd1;
        'd2439 :data = 'd1;
        'd2440 :data = 'd0;
        'd2441 :data = 'd1;
        'd2442 :data = 'd1;
        'd2443 :data = 'd1;
        'd2444 :data = 'd1;
        'd2445 :data = 'd0;
        'd2446 :data = 'd0;
        'd2447 :data = 'd0;
        'd2448 :data = 'd1;
        'd2449 :data = 'd0;
        'd2450 :data = 'd1;
        'd2451 :data = 'd1;
        'd2452 :data = 'd1;
        'd2453 :data = 'd1;
        'd2454 :data = 'd1;
        'd2455 :data = 'd1;
        'd2456 :data = 'd1;
        'd2457 :data = 'd0;
        'd2458 :data = 'd0;
        'd2459 :data = 'd0;
        'd2460 :data = 'd0;
        'd2461 :data = 'd1;
        'd2462 :data = 'd1;
        'd2463 :data = 'd1;
        'd2464 :data = 'd1;
        'd2465 :data = 'd0;
        'd2466 :data = 'd0;
        'd2467 :data = 'd0;
        'd2468 :data = 'd1;
        'd2469 :data = 'd1;
        'd2470 :data = 'd0;
        'd2471 :data = 'd0;
        'd2472 :data = 'd1;
        'd2473 :data = 'd1;
        'd2474 :data = 'd0;
        'd2475 :data = 'd0;
        'd2476 :data = 'd1;
        'd2477 :data = 'd0;
        'd2478 :data = 'd1;
        'd2479 :data = 'd0;
        'd2480 :data = 'd1;
        'd2481 :data = 'd0;
        'd2482 :data = 'd1;
        'd2483 :data = 'd1;
        'd2484 :data = 'd1;
        'd2485 :data = 'd0;
        'd2486 :data = 'd1;
        'd2487 :data = 'd0;
        'd2488 :data = 'd0;
        'd2489 :data = 'd0;
        'd2490 :data = 'd0;
        'd2491 :data = 'd1;
        'd2492 :data = 'd1;
        'd2493 :data = 'd0;
        'd2494 :data = 'd1;
        'd2495 :data = 'd1;
        'd2496 :data = 'd0;
        'd2497 :data = 'd1;
        'd2498 :data = 'd0;
        'd2499 :data = 'd0;
        'd2500 :data = 'd1;
        'd2501 :data = 'd0;
        'd2502 :data = 'd1;
        'd2503 :data = 'd0;
        'd2504 :data = 'd0;
        'd2505 :data = 'd1;
        'd2506 :data = 'd1;
        'd2507 :data = 'd1;
        'd2508 :data = 'd0;
        'd2509 :data = 'd0;
        'd2510 :data = 'd1;
        'd2511 :data = 'd1;
        'd2512 :data = 'd1;
        'd2513 :data = 'd0;
        'd2514 :data = 'd0;
        'd2515 :data = 'd1;
        'd2516 :data = 'd0;
        'd2517 :data = 'd0;
        'd2518 :data = 'd0;
        'd2519 :data = 'd0;
        'd2520 :data = 'd1;
        'd2521 :data = 'd0;
        'd2522 :data = 'd1;
        'd2523 :data = 'd1;
        'd2524 :data = 'd1;
        'd2525 :data = 'd0;
        'd2526 :data = 'd0;
        'd2527 :data = 'd1;
        'd2528 :data = 'd1;
        'd2529 :data = 'd1;
        'd2530 :data = 'd1;
        'd2531 :data = 'd0;
        'd2532 :data = 'd1;
        'd2533 :data = 'd0;
        'd2534 :data = 'd0;
        'd2535 :data = 'd0;
        'd2536 :data = 'd1;
        'd2537 :data = 'd0;
        'd2538 :data = 'd0;
        'd2539 :data = 'd0;
        'd2540 :data = 'd1;
        'd2541 :data = 'd0;
        'd2542 :data = 'd1;
        'd2543 :data = 'd1;
        'd2544 :data = 'd0;
        'd2545 :data = 'd0;
        'd2546 :data = 'd1;
        'd2547 :data = 'd1;
        'd2548 :data = 'd0;
        'd2549 :data = 'd0;
        'd2550 :data = 'd1;
        'd2551 :data = 'd1;
        'd2552 :data = 'd0;
        'd2553 :data = 'd0;
        'd2554 :data = 'd0;
        'd2555 :data = 'd1;
        'd2556 :data = 'd1;
        'd2557 :data = 'd0;
        'd2558 :data = 'd0;
        'd2559 :data = 'd0;
        'd2560 :data = 'd1;
        'd2561 :data = 'd0;
        'd2562 :data = 'd1;
        'd2563 :data = 'd0;
        'd2564 :data = 'd1;
        'd2565 :data = 'd1;
        'd2566 :data = 'd1;
        'd2567 :data = 'd0;
        'd2568 :data = 'd1;
        'd2569 :data = 'd0;
        'd2570 :data = 'd1;
        'd2571 :data = 'd0;
        'd2572 :data = 'd0;
        'd2573 :data = 'd0;
        'd2574 :data = 'd1;
        'd2575 :data = 'd1;
        'd2576 :data = 'd0;
        'd2577 :data = 'd0;
        'd2578 :data = 'd0;
        'd2579 :data = 'd0;
        'd2580 :data = 'd0;
        'd2581 :data = 'd1;
        'd2582 :data = 'd0;
        'd2583 :data = 'd0;
        'd2584 :data = 'd1;
        'd2585 :data = 'd0;
        'd2586 :data = 'd1;
        'd2587 :data = 'd1;
        'd2588 :data = 'd1;
        'd2589 :data = 'd0;
        'd2590 :data = 'd0;
        'd2591 :data = 'd1;
        'd2592 :data = 'd1;
        'd2593 :data = 'd1;
        'd2594 :data = 'd0;
        'd2595 :data = 'd0;
        'd2596 :data = 'd0;
        'd2597 :data = 'd1;
        'd2598 :data = 'd1;
        'd2599 :data = 'd0;
        'd2600 :data = 'd0;
        'd2601 :data = 'd0;
        'd2602 :data = 'd1;
        'd2603 :data = 'd0;
        'd2604 :data = 'd0;
        'd2605 :data = 'd1;
        'd2606 :data = 'd1;
        'd2607 :data = 'd0;
        'd2608 :data = 'd0;
        'd2609 :data = 'd1;
        'd2610 :data = 'd1;
        'd2611 :data = 'd0;
        'd2612 :data = 'd1;
        'd2613 :data = 'd1;
        'd2614 :data = 'd1;
        'd2615 :data = 'd1;
        'd2616 :data = 'd0;
        'd2617 :data = 'd0;
        'd2618 :data = 'd0;
        'd2619 :data = 'd0;
        'd2620 :data = 'd1;
        'd2621 :data = 'd0;
        'd2622 :data = 'd1;
        'd2623 :data = 'd0;
        'd2624 :data = 'd1;
        'd2625 :data = 'd1;
        'd2626 :data = 'd1;
        'd2627 :data = 'd1;
        'd2628 :data = 'd0;
        'd2629 :data = 'd0;
        'd2630 :data = 'd1;
        'd2631 :data = 'd1;
        'd2632 :data = 'd0;
        'd2633 :data = 'd1;
        'd2634 :data = 'd0;
        'd2635 :data = 'd0;
        'd2636 :data = 'd1;
        'd2637 :data = 'd1;
        'd2638 :data = 'd0;
        'd2639 :data = 'd1;
        'd2640 :data = 'd1;
        'd2641 :data = 'd0;
        'd2642 :data = 'd1;
        'd2643 :data = 'd0;
        'd2644 :data = 'd1;
        'd2645 :data = 'd0;
        'd2646 :data = 'd1;
        'd2647 :data = 'd0;
        'd2648 :data = 'd1;
        'd2649 :data = 'd1;
        'd2650 :data = 'd1;
        'd2651 :data = 'd0;
        'd2652 :data = 'd0;
        'd2653 :data = 'd1;
        'd2654 :data = 'd0;
        'd2655 :data = 'd1;
        'd2656 :data = 'd1;
        'd2657 :data = 'd1;
        'd2658 :data = 'd1;
        'd2659 :data = 'd0;
        'd2660 :data = 'd0;
        'd2661 :data = 'd1;
        'd2662 :data = 'd0;
        'd2663 :data = 'd1;
        'd2664 :data = 'd0;
        'd2665 :data = 'd1;
        'd2666 :data = 'd0;
        'd2667 :data = 'd0;
        'd2668 :data = 'd1;
        'd2669 :data = 'd1;
        'd2670 :data = 'd0;
        'd2671 :data = 'd0;
        'd2672 :data = 'd1;
        'd2673 :data = 'd0;
        'd2674 :data = 'd1;
        'd2675 :data = 'd0;
        'd2676 :data = 'd0;
        'd2677 :data = 'd1;
        'd2678 :data = 'd1;
        'd2679 :data = 'd1;
        'd2680 :data = 'd1;
        'd2681 :data = 'd0;
        'd2682 :data = 'd1;
        'd2683 :data = 'd0;
        'd2684 :data = 'd0;
        'd2685 :data = 'd1;
        'd2686 :data = 'd0;
        'd2687 :data = 'd1;
        'd2688 :data = 'd0;
        'd2689 :data = 'd1;
        'd2690 :data = 'd0;
        'd2691 :data = 'd1;
        'd2692 :data = 'd0;
        'd2693 :data = 'd0;
        'd2694 :data = 'd1;
        'd2695 :data = 'd1;
        'd2696 :data = 'd1;
        'd2697 :data = 'd0;
        'd2698 :data = 'd1;
        'd2699 :data = 'd0;
        'd2700 :data = 'd1;
        'd2701 :data = 'd1;
        'd2702 :data = 'd0;
        'd2703 :data = 'd1;
        'd2704 :data = 'd0;
        'd2705 :data = 'd0;
        'd2706 :data = 'd1;
        'd2707 :data = 'd0;
        'd2708 :data = 'd1;
        'd2709 :data = 'd1;
        'd2710 :data = 'd1;
        'd2711 :data = 'd0;
        'd2712 :data = 'd0;
        'd2713 :data = 'd0;
        'd2714 :data = 'd0;
        'd2715 :data = 'd1;
        'd2716 :data = 'd0;
        'd2717 :data = 'd0;
        'd2718 :data = 'd0;
        'd2719 :data = 'd0;
        'd2720 :data = 'd1;
        'd2721 :data = 'd0;
        'd2722 :data = 'd0;
        'd2723 :data = 'd0;
        'd2724 :data = 'd1;
        'd2725 :data = 'd0;
        'd2726 :data = 'd1;
        'd2727 :data = 'd1;
        'd2728 :data = 'd0;
        'd2729 :data = 'd0;
        'd2730 :data = 'd0;
        'd2731 :data = 'd1;
        'd2732 :data = 'd0;
        'd2733 :data = 'd1;
        'd2734 :data = 'd0;
        'd2735 :data = 'd1;
        'd2736 :data = 'd0;
        'd2737 :data = 'd1;
        'd2738 :data = 'd0;
        'd2739 :data = 'd1;
        'd2740 :data = 'd0;
        'd2741 :data = 'd1;
        'd2742 :data = 'd1;
        'd2743 :data = 'd1;
        'd2744 :data = 'd1;
        'd2745 :data = 'd0;
        'd2746 :data = 'd0;
        'd2747 :data = 'd1;
        'd2748 :data = 'd0;
        'd2749 :data = 'd0;
        'd2750 :data = 'd1;
        'd2751 :data = 'd1;
        'd2752 :data = 'd1;
        'd2753 :data = 'd1;
        'd2754 :data = 'd1;
        'd2755 :data = 'd1;
        'd2756 :data = 'd1;
        'd2757 :data = 'd0;
        'd2758 :data = 'd0;
        'd2759 :data = 'd0;
        'd2760 :data = 'd0;
        'd2761 :data = 'd1;
        'd2762 :data = 'd0;
        'd2763 :data = 'd0;
        'd2764 :data = 'd0;
        'd2765 :data = 'd1;
        'd2766 :data = 'd1;
        'd2767 :data = 'd1;
        'd2768 :data = 'd1;
        'd2769 :data = 'd1;
        'd2770 :data = 'd0;
        'd2771 :data = 'd1;
        'd2772 :data = 'd1;
        'd2773 :data = 'd1;
        'd2774 :data = 'd1;
        'd2775 :data = 'd1;
        'd2776 :data = 'd1;
        'd2777 :data = 'd1;
        'd2778 :data = 'd0;
        'd2779 :data = 'd1;
        'd2780 :data = 'd1;
        'd2781 :data = 'd0;
        'd2782 :data = 'd1;
        'd2783 :data = 'd0;
        'd2784 :data = 'd1;
        'd2785 :data = 'd1;
        'd2786 :data = 'd0;
        'd2787 :data = 'd0;
        'd2788 :data = 'd1;
        'd2789 :data = 'd0;
        'd2790 :data = 'd0;
        'd2791 :data = 'd1;
        'd2792 :data = 'd0;
        'd2793 :data = 'd0;
        'd2794 :data = 'd1;
        'd2795 :data = 'd0;
        'd2796 :data = 'd1;
        'd2797 :data = 'd1;
        'd2798 :data = 'd0;
        'd2799 :data = 'd1;
        'd2800 :data = 'd1;
        'd2801 :data = 'd1;
        'd2802 :data = 'd0;
        'd2803 :data = 'd1;
        'd2804 :data = 'd0;
        'd2805 :data = 'd0;
        'd2806 :data = 'd1;
        'd2807 :data = 'd1;
        'd2808 :data = 'd0;
        'd2809 :data = 'd1;
        'd2810 :data = 'd0;
        'd2811 :data = 'd1;
        'd2812 :data = 'd1;
        'd2813 :data = 'd1;
        'd2814 :data = 'd0;
        'd2815 :data = 'd0;
        'd2816 :data = 'd1;
        'd2817 :data = 'd1;
        'd2818 :data = 'd0;
        'd2819 :data = 'd0;
        'd2820 :data = 'd0;
        'd2821 :data = 'd0;
        'd2822 :data = 'd1;
        'd2823 :data = 'd0;
        'd2824 :data = 'd1;
        'd2825 :data = 'd0;
        'd2826 :data = 'd0;
        'd2827 :data = 'd1;
        'd2828 :data = 'd1;
        'd2829 :data = 'd1;
        'd2830 :data = 'd1;
        'd2831 :data = 'd1;
        'd2832 :data = 'd0;
        'd2833 :data = 'd0;
        'd2834 :data = 'd0;
        'd2835 :data = 'd1;
        'd2836 :data = 'd0;
        'd2837 :data = 'd0;
        'd2838 :data = 'd0;
        'd2839 :data = 'd0;
        'd2840 :data = 'd1;
        'd2841 :data = 'd1;
        'd2842 :data = 'd1;
        'd2843 :data = 'd0;
        'd2844 :data = 'd1;
        'd2845 :data = 'd1;
        'd2846 :data = 'd0;
        'd2847 :data = 'd0;
        'd2848 :data = 'd1;
        'd2849 :data = 'd1;
        'd2850 :data = 'd1;
        'd2851 :data = 'd0;
        'd2852 :data = 'd0;
        'd2853 :data = 'd0;
        'd2854 :data = 'd0;
        'd2855 :data = 'd0;
        'd2856 :data = 'd0;
        'd2857 :data = 'd0;
        'd2858 :data = 'd0;
        'd2859 :data = 'd0;
        'd2860 :data = 'd1;
        'd2861 :data = 'd0;
        'd2862 :data = 'd0;
        'd2863 :data = 'd0;
        'd2864 :data = 'd1;
        'd2865 :data = 'd1;
        'd2866 :data = 'd1;
        'd2867 :data = 'd1;
        'd2868 :data = 'd1;
        'd2869 :data = 'd0;
        'd2870 :data = 'd1;
        'd2871 :data = 'd1;
        'd2872 :data = 'd0;
        'd2873 :data = 'd0;
        'd2874 :data = 'd0;
        'd2875 :data = 'd1;
        'd2876 :data = 'd0;
        'd2877 :data = 'd0;
        'd2878 :data = 'd0;
        'd2879 :data = 'd0;
        'd2880 :data = 'd1;
        'd2881 :data = 'd0;
        'd2882 :data = 'd1;
        'd2883 :data = 'd1;
        'd2884 :data = 'd1;
        'd2885 :data = 'd1;
        'd2886 :data = 'd0;
        'd2887 :data = 'd0;
        'd2888 :data = 'd0;
        'd2889 :data = 'd1;
        'd2890 :data = 'd0;
        'd2891 :data = 'd0;
        'd2892 :data = 'd1;
        'd2893 :data = 'd0;
        'd2894 :data = 'd0;
        'd2895 :data = 'd0;
        'd2896 :data = 'd0;
        'd2897 :data = 'd0;
        'd2898 :data = 'd1;
        'd2899 :data = 'd1;
        'd2900 :data = 'd1;
        'd2901 :data = 'd0;
        'd2902 :data = 'd1;
        'd2903 :data = 'd0;
        'd2904 :data = 'd1;
        'd2905 :data = 'd0;
        'd2906 :data = 'd1;
        'd2907 :data = 'd0;
        'd2908 :data = 'd0;
        'd2909 :data = 'd1;
        'd2910 :data = 'd1;
        'd2911 :data = 'd0;
        'd2912 :data = 'd1;
        'd2913 :data = 'd0;
        'd2914 :data = 'd0;
        'd2915 :data = 'd0;
        'd2916 :data = 'd0;
        'd2917 :data = 'd0;
        'd2918 :data = 'd0;
        'd2919 :data = 'd0;
        'd2920 :data = 'd0;
        'd2921 :data = 'd0;
        'd2922 :data = 'd0;
        'd2923 :data = 'd0;
        'd2924 :data = 'd1;
        'd2925 :data = 'd1;
        'd2926 :data = 'd1;
        'd2927 :data = 'd0;
        'd2928 :data = 'd1;
        'd2929 :data = 'd1;
        'd2930 :data = 'd0;
        'd2931 :data = 'd0;
        'd2932 :data = 'd0;
        'd2933 :data = 'd0;
        'd2934 :data = 'd0;
        'd2935 :data = 'd1;
        'd2936 :data = 'd0;
        'd2937 :data = 'd0;
        'd2938 :data = 'd0;
        'd2939 :data = 'd0;
        'd2940 :data = 'd1;
        'd2941 :data = 'd1;
        'd2942 :data = 'd0;
        'd2943 :data = 'd0;
        'd2944 :data = 'd0;
        'd2945 :data = 'd1;
        'd2946 :data = 'd1;
        'd2947 :data = 'd0;
        'd2948 :data = 'd1;
        'd2949 :data = 'd0;
        'd2950 :data = 'd0;
        'd2951 :data = 'd1;
        'd2952 :data = 'd1;
        'd2953 :data = 'd1;
        'd2954 :data = 'd0;
        'd2955 :data = 'd1;
        'd2956 :data = 'd0;
        'd2957 :data = 'd1;
        'd2958 :data = 'd0;
        'd2959 :data = 'd1;
        'd2960 :data = 'd0;
        'd2961 :data = 'd1;
        'd2962 :data = 'd1;
        'd2963 :data = 'd1;
        'd2964 :data = 'd1;
        'd2965 :data = 'd0;
        'd2966 :data = 'd0;
        'd2967 :data = 'd0;
        'd2968 :data = 'd1;
        'd2969 :data = 'd0;
        'd2970 :data = 'd1;
        'd2971 :data = 'd0;
        'd2972 :data = 'd1;
        'd2973 :data = 'd0;
        'd2974 :data = 'd0;
        'd2975 :data = 'd1;
        'd2976 :data = 'd1;
        'd2977 :data = 'd1;
        'd2978 :data = 'd1;
        'd2979 :data = 'd1;
        'd2980 :data = 'd0;
        'd2981 :data = 'd1;
        'd2982 :data = 'd0;
        'd2983 :data = 'd0;
        'd2984 :data = 'd1;
        'd2985 :data = 'd1;
        'd2986 :data = 'd1;
        'd2987 :data = 'd1;
        'd2988 :data = 'd1;
        'd2989 :data = 'd1;
        'd2990 :data = 'd1;
        'd2991 :data = 'd0;
        'd2992 :data = 'd0;
        'd2993 :data = 'd0;
        'd2994 :data = 'd1;
        'd2995 :data = 'd0;
        'd2996 :data = 'd1;
        'd2997 :data = 'd1;
        'd2998 :data = 'd0;
        'd2999 :data = 'd0;
        'd3000 :data = 'd1;
        'd3001 :data = 'd1;
        'd3002 :data = 'd1;
        'd3003 :data = 'd0;
        'd3004 :data = 'd0;
        'd3005 :data = 'd0;
        'd3006 :data = 'd1;
        'd3007 :data = 'd1;
        'd3008 :data = 'd0;
        'd3009 :data = 'd1;
        'd3010 :data = 'd1;
        'd3011 :data = 'd1;
        'd3012 :data = 'd1;
        'd3013 :data = 'd0;
        'd3014 :data = 'd1;
        'd3015 :data = 'd1;
        'd3016 :data = 'd1;
        'd3017 :data = 'd0;
        'd3018 :data = 'd1;
        'd3019 :data = 'd0;
        'd3020 :data = 'd0;
        'd3021 :data = 'd0;
        'd3022 :data = 'd1;
        'd3023 :data = 'd0;
        'd3024 :data = 'd0;
        'd3025 :data = 'd1;
        'd3026 :data = 'd0;
        'd3027 :data = 'd0;
        'd3028 :data = 'd0;
        'd3029 :data = 'd0;
        'd3030 :data = 'd0;
        'd3031 :data = 'd1;
        'd3032 :data = 'd1;
        'd3033 :data = 'd0;
        'd3034 :data = 'd1;
        'd3035 :data = 'd0;
        'd3036 :data = 'd0;
        'd3037 :data = 'd1;
        'd3038 :data = 'd1;
        'd3039 :data = 'd1;
        'd3040 :data = 'd1;
        'd3041 :data = 'd1;
        'd3042 :data = 'd1;
        'd3043 :data = 'd1;
        'd3044 :data = 'd1;
        'd3045 :data = 'd0;
        'd3046 :data = 'd1;
        'd3047 :data = 'd0;
        'd3048 :data = 'd0;
        'd3049 :data = 'd0;
        'd3050 :data = 'd0;
        'd3051 :data = 'd1;
        'd3052 :data = 'd1;
        'd3053 :data = 'd1;
        'd3054 :data = 'd1;
        'd3055 :data = 'd0;
        'd3056 :data = 'd0;
        'd3057 :data = 'd1;
        'd3058 :data = 'd1;
        'd3059 :data = 'd0;
        'd3060 :data = 'd0;
        'd3061 :data = 'd1;
        'd3062 :data = 'd1;
        'd3063 :data = 'd0;
        'd3064 :data = 'd1;
        'd3065 :data = 'd0;
        'd3066 :data = 'd0;
        'd3067 :data = 'd0;
        'd3068 :data = 'd1;
        'd3069 :data = 'd1;
        'd3070 :data = 'd1;
        'd3071 :data = 'd0;
        'd3072 :data = 'd0;
        'd3073 :data = 'd1;
        'd3074 :data = 'd0;
        'd3075 :data = 'd0;
        'd3076 :data = 'd1;
        'd3077 :data = 'd1;
        'd3078 :data = 'd0;
        'd3079 :data = 'd0;
        'd3080 :data = 'd0;
        'd3081 :data = 'd1;
        'd3082 :data = 'd1;
        'd3083 :data = 'd0;
        'd3084 :data = 'd1;
        'd3085 :data = 'd0;
        'd3086 :data = 'd0;
        'd3087 :data = 'd0;
        'd3088 :data = 'd0;
        'd3089 :data = 'd0;
        'd3090 :data = 'd1;
        'd3091 :data = 'd1;
        'd3092 :data = 'd1;
        'd3093 :data = 'd1;
        'd3094 :data = 'd1;
        'd3095 :data = 'd1;
        'd3096 :data = 'd0;
        'd3097 :data = 'd1;
        'd3098 :data = 'd0;
        'd3099 :data = 'd1;
        'd3100 :data = 'd0;
        'd3101 :data = 'd1;
        'd3102 :data = 'd0;
        'd3103 :data = 'd0;
        'd3104 :data = 'd1;
        'd3105 :data = 'd1;
        'd3106 :data = 'd1;
        'd3107 :data = 'd0;
        'd3108 :data = 'd0;
        'd3109 :data = 'd0;
        'd3110 :data = 'd1;
        'd3111 :data = 'd0;
        'd3112 :data = 'd0;
        'd3113 :data = 'd1;
        'd3114 :data = 'd1;
        'd3115 :data = 'd0;
        'd3116 :data = 'd1;
        'd3117 :data = 'd0;
        'd3118 :data = 'd1;
        'd3119 :data = 'd1;
        'd3120 :data = 'd0;
        'd3121 :data = 'd0;
        'd3122 :data = 'd0;
        'd3123 :data = 'd1;
        'd3124 :data = 'd1;
        'd3125 :data = 'd1;
        'd3126 :data = 'd0;
        'd3127 :data = 'd0;
        'd3128 :data = 'd0;
        'd3129 :data = 'd0;
        'd3130 :data = 'd0;
        'd3131 :data = 'd1;
        'd3132 :data = 'd1;
        'd3133 :data = 'd0;
        'd3134 :data = 'd0;
        'd3135 :data = 'd1;
        'd3136 :data = 'd0;
        'd3137 :data = 'd1;
        'd3138 :data = 'd0;
        'd3139 :data = 'd1;
        'd3140 :data = 'd0;
        'd3141 :data = 'd0;
        'd3142 :data = 'd0;
        'd3143 :data = 'd0;
        'd3144 :data = 'd1;
        'd3145 :data = 'd0;
        'd3146 :data = 'd1;
        'd3147 :data = 'd1;
        'd3148 :data = 'd1;
        'd3149 :data = 'd0;
        'd3150 :data = 'd0;
        'd3151 :data = 'd0;
        'd3152 :data = 'd1;
        'd3153 :data = 'd0;
        'd3154 :data = 'd1;
        'd3155 :data = 'd0;
        'd3156 :data = 'd0;
        'd3157 :data = 'd0;
        'd3158 :data = 'd1;
        'd3159 :data = 'd0;
        'd3160 :data = 'd1;
        'd3161 :data = 'd0;
        'd3162 :data = 'd1;
        'd3163 :data = 'd0;
        'd3164 :data = 'd1;
        'd3165 :data = 'd0;
        'd3166 :data = 'd1;
        'd3167 :data = 'd0;
        'd3168 :data = 'd1;
        'd3169 :data = 'd0;
        'd3170 :data = 'd0;
        'd3171 :data = 'd0;
        'd3172 :data = 'd0;
        'd3173 :data = 'd1;
        'd3174 :data = 'd0;
        'd3175 :data = 'd1;
        'd3176 :data = 'd0;
        'd3177 :data = 'd0;
        'd3178 :data = 'd0;
        'd3179 :data = 'd0;
        'd3180 :data = 'd1;
        'd3181 :data = 'd1;
        'd3182 :data = 'd0;
        'd3183 :data = 'd0;
        'd3184 :data = 'd1;
        'd3185 :data = 'd1;
        'd3186 :data = 'd1;
        'd3187 :data = 'd0;
        'd3188 :data = 'd1;
        'd3189 :data = 'd1;
        'd3190 :data = 'd1;
        'd3191 :data = 'd0;
        'd3192 :data = 'd0;
        'd3193 :data = 'd1;
        'd3194 :data = 'd1;
        'd3195 :data = 'd0;
        'd3196 :data = 'd1;
        'd3197 :data = 'd0;
        'd3198 :data = 'd0;
        'd3199 :data = 'd0;
        'd3200 :data = 'd0;
        'd3201 :data = 'd0;
        'd3202 :data = 'd1;
        'd3203 :data = 'd1;
        'd3204 :data = 'd1;
        'd3205 :data = 'd0;
        'd3206 :data = 'd1;
        'd3207 :data = 'd0;
        'd3208 :data = 'd0;
        'd3209 :data = 'd1;
        'd3210 :data = 'd0;
        'd3211 :data = 'd0;
        'd3212 :data = 'd1;
        'd3213 :data = 'd0;
        'd3214 :data = 'd0;
        'd3215 :data = 'd0;
        'd3216 :data = 'd1;
        'd3217 :data = 'd0;
        'd3218 :data = 'd0;
        'd3219 :data = 'd0;
        'd3220 :data = 'd1;
        'd3221 :data = 'd1;
        'd3222 :data = 'd1;
        'd3223 :data = 'd0;
        'd3224 :data = 'd0;
        'd3225 :data = 'd1;
        'd3226 :data = 'd1;
        'd3227 :data = 'd0;
        'd3228 :data = 'd1;
        'd3229 :data = 'd0;
        'd3230 :data = 'd0;
        'd3231 :data = 'd0;
        'd3232 :data = 'd0;
        'd3233 :data = 'd0;
        'd3234 :data = 'd1;
        'd3235 :data = 'd0;
        'd3236 :data = 'd1;
        'd3237 :data = 'd1;
        'd3238 :data = 'd0;
        'd3239 :data = 'd0;
        'd3240 :data = 'd0;
        'd3241 :data = 'd1;
        'd3242 :data = 'd0;
        'd3243 :data = 'd0;
        'd3244 :data = 'd1;
        'd3245 :data = 'd1;
        'd3246 :data = 'd1;
        'd3247 :data = 'd1;
        'd3248 :data = 'd1;
        'd3249 :data = 'd1;
        'd3250 :data = 'd1;
        'd3251 :data = 'd0;
        'd3252 :data = 'd1;
        'd3253 :data = 'd1;
        'd3254 :data = 'd0;
        'd3255 :data = 'd1;
        'd3256 :data = 'd1;
        'd3257 :data = 'd1;
        'd3258 :data = 'd1;
        'd3259 :data = 'd0;
        'd3260 :data = 'd1;
        'd3261 :data = 'd1;
        'd3262 :data = 'd1;
        'd3263 :data = 'd0;
        'd3264 :data = 'd1;
        'd3265 :data = 'd0;
        'd3266 :data = 'd1;
        'd3267 :data = 'd1;
        'd3268 :data = 'd0;
        'd3269 :data = 'd0;
        'd3270 :data = 'd1;
        'd3271 :data = 'd1;
        'd3272 :data = 'd1;
        'd3273 :data = 'd1;
        'd3274 :data = 'd1;
        'd3275 :data = 'd1;
        'd3276 :data = 'd1;
        'd3277 :data = 'd0;
        'd3278 :data = 'd0;
        'd3279 :data = 'd0;
        'd3280 :data = 'd0;
        'd3281 :data = 'd1;
        'd3282 :data = 'd1;
        'd3283 :data = 'd0;
        'd3284 :data = 'd0;
        'd3285 :data = 'd0;
        'd3286 :data = 'd1;
        'd3287 :data = 'd0;
        'd3288 :data = 'd1;
        'd3289 :data = 'd0;
        'd3290 :data = 'd0;
        'd3291 :data = 'd1;
        'd3292 :data = 'd0;
        'd3293 :data = 'd1;
        'd3294 :data = 'd1;
        'd3295 :data = 'd0;
        'd3296 :data = 'd0;
        'd3297 :data = 'd0;
        'd3298 :data = 'd1;
        'd3299 :data = 'd0;
        'd3300 :data = 'd1;
        'd3301 :data = 'd1;
        'd3302 :data = 'd1;
        'd3303 :data = 'd0;
        'd3304 :data = 'd1;
        'd3305 :data = 'd1;
        'd3306 :data = 'd0;
        'd3307 :data = 'd1;
        'd3308 :data = 'd0;
        'd3309 :data = 'd0;
        'd3310 :data = 'd1;
        'd3311 :data = 'd0;
        'd3312 :data = 'd1;
        'd3313 :data = 'd0;
        'd3314 :data = 'd1;
        'd3315 :data = 'd1;
        'd3316 :data = 'd1;
        'd3317 :data = 'd0;
        'd3318 :data = 'd1;
        'd3319 :data = 'd1;
        'd3320 :data = 'd0;
        'd3321 :data = 'd0;
        'd3322 :data = 'd1;
        'd3323 :data = 'd0;
        'd3324 :data = 'd0;
        'd3325 :data = 'd1;
        'd3326 :data = 'd1;
        'd3327 :data = 'd1;
        'd3328 :data = 'd0;
        'd3329 :data = 'd1;
        'd3330 :data = 'd0;
        'd3331 :data = 'd1;
        'd3332 :data = 'd0;
        'd3333 :data = 'd0;
        'd3334 :data = 'd1;
        'd3335 :data = 'd1;
        'd3336 :data = 'd1;
        'd3337 :data = 'd1;
        'd3338 :data = 'd1;
        'd3339 :data = 'd1;
        'd3340 :data = 'd1;
        'd3341 :data = 'd1;
        'd3342 :data = 'd0;
        'd3343 :data = 'd1;
        'd3344 :data = 'd1;
        'd3345 :data = 'd0;
        'd3346 :data = 'd0;
        'd3347 :data = 'd0;
        'd3348 :data = 'd0;
        'd3349 :data = 'd1;
        'd3350 :data = 'd1;
        'd3351 :data = 'd1;
        'd3352 :data = 'd1;
        'd3353 :data = 'd0;
        'd3354 :data = 'd1;
        'd3355 :data = 'd0;
        'd3356 :data = 'd1;
        'd3357 :data = 'd0;
        'd3358 :data = 'd1;
        'd3359 :data = 'd1;
        'd3360 :data = 'd1;
        'd3361 :data = 'd1;
        'd3362 :data = 'd1;
        'd3363 :data = 'd1;
        'd3364 :data = 'd1;
        'd3365 :data = 'd1;
        'd3366 :data = 'd0;
        'd3367 :data = 'd1;
        'd3368 :data = 'd1;
        'd3369 :data = 'd1;
        'd3370 :data = 'd1;
        'd3371 :data = 'd0;
        'd3372 :data = 'd0;
        'd3373 :data = 'd1;
        'd3374 :data = 'd1;
        'd3375 :data = 'd0;
        'd3376 :data = 'd0;
        'd3377 :data = 'd0;
        'd3378 :data = 'd0;
        'd3379 :data = 'd0;
        'd3380 :data = 'd0;
        'd3381 :data = 'd1;
        'd3382 :data = 'd0;
        'd3383 :data = 'd0;
        'd3384 :data = 'd0;
        'd3385 :data = 'd0;
        'd3386 :data = 'd1;
        'd3387 :data = 'd1;
        'd3388 :data = 'd1;
        'd3389 :data = 'd1;
        'd3390 :data = 'd1;
        'd3391 :data = 'd0;
        'd3392 :data = 'd0;
        'd3393 :data = 'd1;
        'd3394 :data = 'd0;
        'd3395 :data = 'd0;
        'd3396 :data = 'd0;
        'd3397 :data = 'd0;
        'd3398 :data = 'd1;
        'd3399 :data = 'd1;
        'd3400 :data = 'd1;
        'd3401 :data = 'd1;
        'd3402 :data = 'd1;
        'd3403 :data = 'd0;
        'd3404 :data = 'd0;
        'd3405 :data = 'd1;
        'd3406 :data = 'd0;
        'd3407 :data = 'd0;
        'd3408 :data = 'd0;
        'd3409 :data = 'd1;
        'd3410 :data = 'd0;
        'd3411 :data = 'd1;
        'd3412 :data = 'd0;
        'd3413 :data = 'd0;
        'd3414 :data = 'd1;
        'd3415 :data = 'd0;
        'd3416 :data = 'd1;
        'd3417 :data = 'd0;
        'd3418 :data = 'd1;
        'd3419 :data = 'd1;
        'd3420 :data = 'd1;
        'd3421 :data = 'd1;
        'd3422 :data = 'd0;
        'd3423 :data = 'd1;
        'd3424 :data = 'd0;
        'd3425 :data = 'd0;
        'd3426 :data = 'd0;
        'd3427 :data = 'd1;
        'd3428 :data = 'd1;
        'd3429 :data = 'd1;
        'd3430 :data = 'd0;
        'd3431 :data = 'd1;
        'd3432 :data = 'd0;
        'd3433 :data = 'd0;
        'd3434 :data = 'd1;
        'd3435 :data = 'd1;
        'd3436 :data = 'd0;
        'd3437 :data = 'd1;
        'd3438 :data = 'd0;
        'd3439 :data = 'd1;
        'd3440 :data = 'd0;
        'd3441 :data = 'd1;
        'd3442 :data = 'd0;
        'd3443 :data = 'd0;
        'd3444 :data = 'd1;
        'd3445 :data = 'd0;
        'd3446 :data = 'd0;
        'd3447 :data = 'd1;
        'd3448 :data = 'd1;
        'd3449 :data = 'd1;
        'd3450 :data = 'd0;
        'd3451 :data = 'd1;
        'd3452 :data = 'd0;
        'd3453 :data = 'd0;
        'd3454 :data = 'd0;
        'd3455 :data = 'd1;
        'd3456 :data = 'd1;
        'd3457 :data = 'd0;
        'd3458 :data = 'd1;
        'd3459 :data = 'd1;
        'd3460 :data = 'd1;
        'd3461 :data = 'd1;
        'd3462 :data = 'd0;
        'd3463 :data = 'd0;
        'd3464 :data = 'd0;
        'd3465 :data = 'd0;
        'd3466 :data = 'd0;
        'd3467 :data = 'd1;
        'd3468 :data = 'd0;
        'd3469 :data = 'd0;
        'd3470 :data = 'd1;
        'd3471 :data = 'd0;
        'd3472 :data = 'd0;
        'd3473 :data = 'd1;
        'd3474 :data = 'd0;
        'd3475 :data = 'd0;
        'd3476 :data = 'd0;
        'd3477 :data = 'd1;
        'd3478 :data = 'd0;
        'd3479 :data = 'd0;
        'd3480 :data = 'd0;
        'd3481 :data = 'd1;
        'd3482 :data = 'd1;
        'd3483 :data = 'd0;
        'd3484 :data = 'd1;
        'd3485 :data = 'd1;
        'd3486 :data = 'd0;
        'd3487 :data = 'd1;
        'd3488 :data = 'd0;
        'd3489 :data = 'd0;
        'd3490 :data = 'd0;
        'd3491 :data = 'd1;
        'd3492 :data = 'd0;
        'd3493 :data = 'd1;
        'd3494 :data = 'd1;
        'd3495 :data = 'd1;
        'd3496 :data = 'd0;
        'd3497 :data = 'd0;
        'd3498 :data = 'd0;
        'd3499 :data = 'd1;
        'd3500 :data = 'd1;
        'd3501 :data = 'd1;
        'd3502 :data = 'd1;
        'd3503 :data = 'd0;
        'd3504 :data = 'd0;
        'd3505 :data = 'd1;
        'd3506 :data = 'd1;
        'd3507 :data = 'd1;
        'd3508 :data = 'd0;
        'd3509 :data = 'd1;
        'd3510 :data = 'd0;
        'd3511 :data = 'd1;
        'd3512 :data = 'd1;
        'd3513 :data = 'd1;
        'd3514 :data = 'd0;
        'd3515 :data = 'd1;
        'd3516 :data = 'd1;
        'd3517 :data = 'd1;
        'd3518 :data = 'd0;
        'd3519 :data = 'd0;
        'd3520 :data = 'd1;
        'd3521 :data = 'd1;
        'd3522 :data = 'd1;
        'd3523 :data = 'd0;
        'd3524 :data = 'd1;
        'd3525 :data = 'd1;
        'd3526 :data = 'd1;
        'd3527 :data = 'd0;
        'd3528 :data = 'd1;
        'd3529 :data = 'd1;
        'd3530 :data = 'd1;
        'd3531 :data = 'd0;
        'd3532 :data = 'd1;
        'd3533 :data = 'd0;
        'd3534 :data = 'd1;
        'd3535 :data = 'd0;
        'd3536 :data = 'd1;
        'd3537 :data = 'd0;
        'd3538 :data = 'd0;
        'd3539 :data = 'd0;
        'd3540 :data = 'd1;
        'd3541 :data = 'd0;
        'd3542 :data = 'd0;
        'd3543 :data = 'd1;
        'd3544 :data = 'd1;
        'd3545 :data = 'd0;
        'd3546 :data = 'd1;
        'd3547 :data = 'd0;
        'd3548 :data = 'd0;
        'd3549 :data = 'd0;
        'd3550 :data = 'd1;
        'd3551 :data = 'd0;
        'd3552 :data = 'd0;
        'd3553 :data = 'd1;
        'd3554 :data = 'd0;
        'd3555 :data = 'd0;
        'd3556 :data = 'd0;
        'd3557 :data = 'd0;
        'd3558 :data = 'd1;
        'd3559 :data = 'd0;
        'd3560 :data = 'd0;
        'd3561 :data = 'd1;
        'd3562 :data = 'd1;
        'd3563 :data = 'd0;
        'd3564 :data = 'd0;
        'd3565 :data = 'd1;
        'd3566 :data = 'd0;
        'd3567 :data = 'd1;
        'd3568 :data = 'd1;
        'd3569 :data = 'd1;
        'd3570 :data = 'd0;
        'd3571 :data = 'd0;
        'd3572 :data = 'd1;
        'd3573 :data = 'd1;
        'd3574 :data = 'd1;
        'd3575 :data = 'd0;
        'd3576 :data = 'd0;
        'd3577 :data = 'd0;
        'd3578 :data = 'd0;
        'd3579 :data = 'd1;
        'd3580 :data = 'd0;
        'd3581 :data = 'd0;
        'd3582 :data = 'd1;
        'd3583 :data = 'd1;
        'd3584 :data = 'd0;
        'd3585 :data = 'd0;
        'd3586 :data = 'd0;
        'd3587 :data = 'd1;
        'd3588 :data = 'd0;
        'd3589 :data = 'd0;
        'd3590 :data = 'd1;
        'd3591 :data = 'd1;
        'd3592 :data = 'd1;
        'd3593 :data = 'd0;
        'd3594 :data = 'd0;
        'd3595 :data = 'd1;
        'd3596 :data = 'd0;
        'd3597 :data = 'd1;
        'd3598 :data = 'd1;
        'd3599 :data = 'd0;
        'd3600 :data = 'd1;
        'd3601 :data = 'd0;
        'd3602 :data = 'd0;
        'd3603 :data = 'd0;
        'd3604 :data = 'd0;
        'd3605 :data = 'd1;
        'd3606 :data = 'd0;
        'd3607 :data = 'd1;
        'd3608 :data = 'd0;
        'd3609 :data = 'd1;
        'd3610 :data = 'd1;
        'd3611 :data = 'd1;
        'd3612 :data = 'd1;
        'd3613 :data = 'd1;
        'd3614 :data = 'd1;
        'd3615 :data = 'd1;
        'd3616 :data = 'd0;
        'd3617 :data = 'd1;
        'd3618 :data = 'd1;
        'd3619 :data = 'd1;
        'd3620 :data = 'd0;
        'd3621 :data = 'd1;
        'd3622 :data = 'd1;
        'd3623 :data = 'd0;
        'd3624 :data = 'd0;
        'd3625 :data = 'd1;
        'd3626 :data = 'd0;
        'd3627 :data = 'd1;
        'd3628 :data = 'd0;
        'd3629 :data = 'd0;
        'd3630 :data = 'd1;
        'd3631 :data = 'd0;
        'd3632 :data = 'd1;
        'd3633 :data = 'd1;
        'd3634 :data = 'd1;
        'd3635 :data = 'd0;
        'd3636 :data = 'd1;
        'd3637 :data = 'd0;
        'd3638 :data = 'd0;
        'd3639 :data = 'd1;
        'd3640 :data = 'd0;
        'd3641 :data = 'd1;
        'd3642 :data = 'd1;
        'd3643 :data = 'd0;
        'd3644 :data = 'd0;
        'd3645 :data = 'd1;
        'd3646 :data = 'd0;
        'd3647 :data = 'd0;
        'd3648 :data = 'd1;
        'd3649 :data = 'd1;
        'd3650 :data = 'd0;
        'd3651 :data = 'd0;
        'd3652 :data = 'd0;
        'd3653 :data = 'd1;
        'd3654 :data = 'd1;
        'd3655 :data = 'd0;
        'd3656 :data = 'd0;
        'd3657 :data = 'd0;
        'd3658 :data = 'd0;
        'd3659 :data = 'd0;
        'd3660 :data = 'd0;
        'd3661 :data = 'd0;
        'd3662 :data = 'd0;
        'd3663 :data = 'd1;
        'd3664 :data = 'd1;
        'd3665 :data = 'd1;
        'd3666 :data = 'd0;
        'd3667 :data = 'd0;
        'd3668 :data = 'd1;
        'd3669 :data = 'd1;
        'd3670 :data = 'd0;
        'd3671 :data = 'd0;
        'd3672 :data = 'd1;
        'd3673 :data = 'd0;
        'd3674 :data = 'd1;
        'd3675 :data = 'd1;
        'd3676 :data = 'd0;
        'd3677 :data = 'd1;
        'd3678 :data = 'd0;
        'd3679 :data = 'd0;
        'd3680 :data = 'd0;
        'd3681 :data = 'd1;
        'd3682 :data = 'd0;
        'd3683 :data = 'd1;
        'd3684 :data = 'd1;
        'd3685 :data = 'd1;
        'd3686 :data = 'd0;
        'd3687 :data = 'd1;
        'd3688 :data = 'd1;
        'd3689 :data = 'd1;
        'd3690 :data = 'd0;
        'd3691 :data = 'd0;
        'd3692 :data = 'd0;
        'd3693 :data = 'd1;
        'd3694 :data = 'd1;
        'd3695 :data = 'd1;
        'd3696 :data = 'd1;
        'd3697 :data = 'd1;
        'd3698 :data = 'd1;
        'd3699 :data = 'd1;
        'd3700 :data = 'd0;
        'd3701 :data = 'd1;
        'd3702 :data = 'd0;
        'd3703 :data = 'd1;
        'd3704 :data = 'd0;
        'd3705 :data = 'd1;
        'd3706 :data = 'd1;
        'd3707 :data = 'd0;
        'd3708 :data = 'd1;
        'd3709 :data = 'd0;
        'd3710 :data = 'd0;
        'd3711 :data = 'd1;
        'd3712 :data = 'd1;
        'd3713 :data = 'd1;
        'd3714 :data = 'd1;
        'd3715 :data = 'd1;
        'd3716 :data = 'd1;
        'd3717 :data = 'd0;
        'd3718 :data = 'd0;
        'd3719 :data = 'd0;
        'd3720 :data = 'd1;
        'd3721 :data = 'd0;
        'd3722 :data = 'd0;
        'd3723 :data = 'd0;
        'd3724 :data = 'd1;
        'd3725 :data = 'd0;
        'd3726 :data = 'd0;
        'd3727 :data = 'd0;
        'd3728 :data = 'd1;
        'd3729 :data = 'd1;
        'd3730 :data = 'd0;
        'd3731 :data = 'd1;
        'd3732 :data = 'd0;
        'd3733 :data = 'd1;
        'd3734 :data = 'd1;
        'd3735 :data = 'd0;
        'd3736 :data = 'd1;
        'd3737 :data = 'd1;
        'd3738 :data = 'd1;
        'd3739 :data = 'd0;
        'd3740 :data = 'd1;
        'd3741 :data = 'd1;
        'd3742 :data = 'd0;
        'd3743 :data = 'd1;
        'd3744 :data = 'd0;
        'd3745 :data = 'd1;
        'd3746 :data = 'd0;
        'd3747 :data = 'd0;
        'd3748 :data = 'd1;
        'd3749 :data = 'd1;
        'd3750 :data = 'd1;
        'd3751 :data = 'd0;
        'd3752 :data = 'd1;
        'd3753 :data = 'd0;
        'd3754 :data = 'd0;
        'd3755 :data = 'd0;
        'd3756 :data = 'd0;
        'd3757 :data = 'd1;
        'd3758 :data = 'd0;
        'd3759 :data = 'd0;
        'd3760 :data = 'd0;
        'd3761 :data = 'd1;
        'd3762 :data = 'd0;
        'd3763 :data = 'd0;
        'd3764 :data = 'd0;
        'd3765 :data = 'd1;
        'd3766 :data = 'd1;
        'd3767 :data = 'd1;
        'd3768 :data = 'd0;
        'd3769 :data = 'd1;
        'd3770 :data = 'd1;
        'd3771 :data = 'd1;
        'd3772 :data = 'd1;
        'd3773 :data = 'd0;
        'd3774 :data = 'd1;
        'd3775 :data = 'd1;
        'd3776 :data = 'd1;
        'd3777 :data = 'd1;
        'd3778 :data = 'd1;
        'd3779 :data = 'd0;
        'd3780 :data = 'd1;
        'd3781 :data = 'd0;
        'd3782 :data = 'd0;
        'd3783 :data = 'd0;
        'd3784 :data = 'd0;
        'd3785 :data = 'd0;
        'd3786 :data = 'd1;
        'd3787 :data = 'd0;
        'd3788 :data = 'd0;
        'd3789 :data = 'd1;
        'd3790 :data = 'd0;
        'd3791 :data = 'd1;
        'd3792 :data = 'd0;
        'd3793 :data = 'd0;
        'd3794 :data = 'd0;
        'd3795 :data = 'd0;
        'd3796 :data = 'd0;
        'd3797 :data = 'd0;
        'd3798 :data = 'd1;
        'd3799 :data = 'd0;
        'd3800 :data = 'd0;
        'd3801 :data = 'd0;
        'd3802 :data = 'd1;
        'd3803 :data = 'd1;
        'd3804 :data = 'd0;
        'd3805 :data = 'd1;
        'd3806 :data = 'd0;
        'd3807 :data = 'd1;
        'd3808 :data = 'd1;
        'd3809 :data = 'd1;
        'd3810 :data = 'd1;
        'd3811 :data = 'd1;
        'd3812 :data = 'd1;
        'd3813 :data = 'd1;
        'd3814 :data = 'd0;
        'd3815 :data = 'd0;
        'd3816 :data = 'd1;
        'd3817 :data = 'd0;
        'd3818 :data = 'd1;
        'd3819 :data = 'd0;
        'd3820 :data = 'd1;
        'd3821 :data = 'd0;
        'd3822 :data = 'd1;
        'd3823 :data = 'd1;
        'd3824 :data = 'd1;
        'd3825 :data = 'd1;
        'd3826 :data = 'd1;
        'd3827 :data = 'd0;
        'd3828 :data = 'd0;
        'd3829 :data = 'd0;
        'd3830 :data = 'd1;
        'd3831 :data = 'd0;
        'd3832 :data = 'd1;
        'd3833 :data = 'd1;
        'd3834 :data = 'd1;
        'd3835 :data = 'd1;
        'd3836 :data = 'd1;
        'd3837 :data = 'd1;
        'd3838 :data = 'd0;
        'd3839 :data = 'd0;
        'd3840 :data = 'd1;
        'd3841 :data = 'd0;
        'd3842 :data = 'd1;
        'd3843 :data = 'd1;
        'd3844 :data = 'd0;
        'd3845 :data = 'd1;
        'd3846 :data = 'd0;
        'd3847 :data = 'd0;
        'd3848 :data = 'd1;
        'd3849 :data = 'd1;
        'd3850 :data = 'd0;
        'd3851 :data = 'd1;
        'd3852 :data = 'd1;
        'd3853 :data = 'd0;
        'd3854 :data = 'd0;
        'd3855 :data = 'd0;
        'd3856 :data = 'd1;
        'd3857 :data = 'd0;
        'd3858 :data = 'd1;
        'd3859 :data = 'd0;
        'd3860 :data = 'd1;
        'd3861 :data = 'd0;
        'd3862 :data = 'd0;
        'd3863 :data = 'd0;
        'd3864 :data = 'd1;
        'd3865 :data = 'd0;
        'd3866 :data = 'd1;
        'd3867 :data = 'd1;
        'd3868 :data = 'd0;
        'd3869 :data = 'd1;
        'd3870 :data = 'd1;
        'd3871 :data = 'd0;
        'd3872 :data = 'd0;
        'd3873 :data = 'd1;
        'd3874 :data = 'd0;
        'd3875 :data = 'd1;
        'd3876 :data = 'd0;
        'd3877 :data = 'd1;
        'd3878 :data = 'd0;
        'd3879 :data = 'd0;
        'd3880 :data = 'd1;
        'd3881 :data = 'd0;
        'd3882 :data = 'd1;
        'd3883 :data = 'd0;
        'd3884 :data = 'd0;
        'd3885 :data = 'd0;
        'd3886 :data = 'd0;
        'd3887 :data = 'd1;
        'd3888 :data = 'd1;
        'd3889 :data = 'd1;
        'd3890 :data = 'd0;
        'd3891 :data = 'd0;
        'd3892 :data = 'd1;
        'd3893 :data = 'd0;
        'd3894 :data = 'd0;
        'd3895 :data = 'd0;
        'd3896 :data = 'd1;
        'd3897 :data = 'd0;
        'd3898 :data = 'd0;
        'd3899 :data = 'd1;
        'd3900 :data = 'd1;
        'd3901 :data = 'd0;
        'd3902 :data = 'd1;
        'd3903 :data = 'd1;
        'd3904 :data = 'd1;
        'd3905 :data = 'd0;
        'd3906 :data = 'd1;
        'd3907 :data = 'd1;
        'd3908 :data = 'd1;
        'd3909 :data = 'd1;
        'd3910 :data = 'd0;
        'd3911 :data = 'd0;
        'd3912 :data = 'd0;
        'd3913 :data = 'd1;
        'd3914 :data = 'd1;
        'd3915 :data = 'd1;
        'd3916 :data = 'd1;
        'd3917 :data = 'd1;
        'd3918 :data = 'd0;
        'd3919 :data = 'd0;
        'd3920 :data = 'd0;
        'd3921 :data = 'd0;
        'd3922 :data = 'd1;
        'd3923 :data = 'd1;
        'd3924 :data = 'd1;
        'd3925 :data = 'd1;
        'd3926 :data = 'd0;
        'd3927 :data = 'd0;
        'd3928 :data = 'd0;
        'd3929 :data = 'd0;
        'd3930 :data = 'd1;
        'd3931 :data = 'd0;
        'd3932 :data = 'd1;
        'd3933 :data = 'd1;
        'd3934 :data = 'd1;
        'd3935 :data = 'd1;
        'd3936 :data = 'd0;
        'd3937 :data = 'd0;
        'd3938 :data = 'd1;
        'd3939 :data = 'd1;
        'd3940 :data = 'd0;
        'd3941 :data = 'd0;
        'd3942 :data = 'd1;
        'd3943 :data = 'd1;
        'd3944 :data = 'd0;
        'd3945 :data = 'd1;
        'd3946 :data = 'd0;
        'd3947 :data = 'd0;
        'd3948 :data = 'd0;
        'd3949 :data = 'd1;
        'd3950 :data = 'd1;
        'd3951 :data = 'd0;
        'd3952 :data = 'd1;
        'd3953 :data = 'd1;
        'd3954 :data = 'd0;
        'd3955 :data = 'd0;
        'd3956 :data = 'd0;
        'd3957 :data = 'd1;
        'd3958 :data = 'd1;
        'd3959 :data = 'd0;
        'd3960 :data = 'd1;
        'd3961 :data = 'd0;
        'd3962 :data = 'd0;
        'd3963 :data = 'd1;
        'd3964 :data = 'd1;
        'd3965 :data = 'd1;
        'd3966 :data = 'd1;
        'd3967 :data = 'd0;
        'd3968 :data = 'd0;
        'd3969 :data = 'd1;
        'd3970 :data = 'd1;
        'd3971 :data = 'd1;
        'd3972 :data = 'd1;
        'd3973 :data = 'd0;
        'd3974 :data = 'd1;
        'd3975 :data = 'd1;
        'd3976 :data = 'd0;
        'd3977 :data = 'd1;
        'd3978 :data = 'd0;
        'd3979 :data = 'd1;
        'd3980 :data = 'd0;
        'd3981 :data = 'd1;
        'd3982 :data = 'd0;
        'd3983 :data = 'd1;
        'd3984 :data = 'd1;
        'd3985 :data = 'd1;
        'd3986 :data = 'd1;
        'd3987 :data = 'd1;
        'd3988 :data = 'd1;
        'd3989 :data = 'd1;
        'd3990 :data = 'd0;
        'd3991 :data = 'd0;
        'd3992 :data = 'd0;
        'd3993 :data = 'd1;
        'd3994 :data = 'd1;
        'd3995 :data = 'd1;
        'd3996 :data = 'd1;
        'd3997 :data = 'd0;
        'd3998 :data = 'd1;
        'd3999 :data = 'd0;
        'd4000 :data = 'd1;
        'd4001 :data = 'd0;
        'd4002 :data = 'd1;
        'd4003 :data = 'd1;
        'd4004 :data = 'd1;
        'd4005 :data = 'd1;
        'd4006 :data = 'd1;
        'd4007 :data = 'd0;
        'd4008 :data = 'd1;
        'd4009 :data = 'd0;
        'd4010 :data = 'd0;
        'd4011 :data = 'd0;
        'd4012 :data = 'd1;
        'd4013 :data = 'd0;
        'd4014 :data = 'd1;
        'd4015 :data = 'd1;
        'd4016 :data = 'd0;
        'd4017 :data = 'd1;
        'd4018 :data = 'd0;
        'd4019 :data = 'd0;
        'd4020 :data = 'd0;
        'd4021 :data = 'd1;
        'd4022 :data = 'd1;
        'd4023 :data = 'd1;
        'd4024 :data = 'd1;
        'd4025 :data = 'd1;
        'd4026 :data = 'd1;
        'd4027 :data = 'd1;
        'd4028 :data = 'd1;
        'd4029 :data = 'd0;
        'd4030 :data = 'd1;
        'd4031 :data = 'd1;
        'd4032 :data = 'd0;
        'd4033 :data = 'd1;
        'd4034 :data = 'd0;
        'd4035 :data = 'd1;
        'd4036 :data = 'd1;
        'd4037 :data = 'd1;
        'd4038 :data = 'd1;
        'd4039 :data = 'd1;
        'd4040 :data = 'd1;
        'd4041 :data = 'd1;
        'd4042 :data = 'd0;
        'd4043 :data = 'd1;
        'd4044 :data = 'd0;
        'd4045 :data = 'd1;
        'd4046 :data = 'd0;
        'd4047 :data = 'd1;
        'd4048 :data = 'd0;
        'd4049 :data = 'd0;
        'd4050 :data = 'd0;
        'd4051 :data = 'd1;
        'd4052 :data = 'd0;
        'd4053 :data = 'd1;
        'd4054 :data = 'd0;
        'd4055 :data = 'd1;
        'd4056 :data = 'd0;
        'd4057 :data = 'd1;
        'd4058 :data = 'd0;
        'd4059 :data = 'd1;
        'd4060 :data = 'd0;
        'd4061 :data = 'd1;
        'd4062 :data = 'd0;
        'd4063 :data = 'd1;
        'd4064 :data = 'd1;
        'd4065 :data = 'd1;
        'd4066 :data = 'd0;
        'd4067 :data = 'd0;
        'd4068 :data = 'd1;
        'd4069 :data = 'd1;
        'd4070 :data = 'd1;
        'd4071 :data = 'd1;
        'd4072 :data = 'd1;
        'd4073 :data = 'd0;
        'd4074 :data = 'd1;
        'd4075 :data = 'd0;
        'd4076 :data = 'd0;
        'd4077 :data = 'd1;
        'd4078 :data = 'd0;
        'd4079 :data = 'd0;
        'd4080 :data = 'd0;
        'd4081 :data = 'd1;
        'd4082 :data = 'd0;
        'd4083 :data = 'd1;
        'd4084 :data = 'd1;
        'd4085 :data = 'd0;
        'd4086 :data = 'd0;
        'd4087 :data = 'd0;
        'd4088 :data = 'd1;
        'd4089 :data = 'd0;
        'd4090 :data = 'd0;
        'd4091 :data = 'd1;
        'd4092 :data = 'd1;
        'd4093 :data = 'd0;
        'd4094 :data = 'd1;
        'd4095 :data = 'd1;
        default: data = 'd0;
    endcase
end
endmodule
