`timescale 1ns/100ps

module pn_rom ( 
// write input and output here
    input               clk,
    input               rst_n,
    input               ena,
    input       [9:0]  address_in,
    output  reg [0:0]  data_out,
    output  reg         valid_out
);

// declare wires and regsiters here
reg [0:0]  data;

// rom table here
always @(posedge clk) begin 
    if (!rst_n) begin
        data_out <= 'b0;
        valid_out <= 'b0;
    end
    else if (!ena) begin
        data_out <= 'b0;
        valid_out <= 'b0;
    end
    else begin
        data_out <= data;
        valid_out <= 1'b1;
    end
end

always @(posedge clk) begin
    case(address_in)
        10'd0 :data = 'b1;
        10'd1 :data = 'b0;
        10'd2 :data = 'b0;
        10'd3 :data = 'b0;
        10'd4 :data = 'b1;
        10'd5 :data = 'b1;
        10'd6 :data = 'b1;
        10'd7 :data = 'b1;
        10'd8 :data = 'b1;
        10'd9 :data = 'b1;
        10'd10 :data = 'b1;
        10'd11 :data = 'b1;
        10'd12 :data = 'b0;
        10'd13 :data = 'b0;
        10'd14 :data = 'b0;
        10'd15 :data = 'b1;
        10'd16 :data = 'b1;
        10'd17 :data = 'b1;
        10'd18 :data = 'b1;
        10'd19 :data = 'b1;
        10'd20 :data = 'b1;
        10'd21 :data = 'b1;
        10'd22 :data = 'b0;
        10'd23 :data = 'b0;
        10'd24 :data = 'b0;
        10'd25 :data = 'b1;
        10'd26 :data = 'b1;
        10'd27 :data = 'b1;
        10'd28 :data = 'b1;
        10'd29 :data = 'b0;
        10'd30 :data = 'b0;
        10'd31 :data = 'b1;
        10'd32 :data = 'b1;
        10'd33 :data = 'b0;
        10'd34 :data = 'b0;
        10'd35 :data = 'b1;
        10'd36 :data = 'b1;
        10'd37 :data = 'b0;
        10'd38 :data = 'b1;
        10'd39 :data = 'b1;
        10'd40 :data = 'b1;
        10'd41 :data = 'b1;
        10'd42 :data = 'b1;
        10'd43 :data = 'b0;
        10'd44 :data = 'b0;
        10'd45 :data = 'b0;
        10'd46 :data = 'b0;
        10'd47 :data = 'b0;
        10'd48 :data = 'b1;
        10'd49 :data = 'b0;
        10'd50 :data = 'b1;
        10'd51 :data = 'b0;
        10'd52 :data = 'b1;
        10'd53 :data = 'b1;
        10'd54 :data = 'b1;
        10'd55 :data = 'b0;
        10'd56 :data = 'b0;
        10'd57 :data = 'b0;
        10'd58 :data = 'b1;
        10'd59 :data = 'b1;
        10'd60 :data = 'b0;
        10'd61 :data = 'b0;
        10'd62 :data = 'b1;
        10'd63 :data = 'b0;
        10'd64 :data = 'b0;
        10'd65 :data = 'b1;
        10'd66 :data = 'b1;
        10'd67 :data = 'b1;
        10'd68 :data = 'b1;
        10'd69 :data = 'b1;
        10'd70 :data = 'b1;
        10'd71 :data = 'b0;
        10'd72 :data = 'b0;
        10'd73 :data = 'b1;
        10'd74 :data = 'b1;
        10'd75 :data = 'b0;
        10'd76 :data = 'b0;
        10'd77 :data = 'b1;
        10'd78 :data = 'b0;
        10'd79 :data = 'b1;
        10'd80 :data = 'b1;
        10'd81 :data = 'b1;
        10'd82 :data = 'b0;
        10'd83 :data = 'b1;
        10'd84 :data = 'b0;
        10'd85 :data = 'b0;
        10'd86 :data = 'b0;
        10'd87 :data = 'b0;
        10'd88 :data = 'b1;
        10'd89 :data = 'b0;
        10'd90 :data = 'b1;
        10'd91 :data = 'b1;
        10'd92 :data = 'b1;
        10'd93 :data = 'b1;
        10'd94 :data = 'b0;
        10'd95 :data = 'b1;
        10'd96 :data = 'b0;
        10'd97 :data = 'b1;
        10'd98 :data = 'b1;
        10'd99 :data = 'b0;
        10'd100 :data = 'b0;
        10'd101 :data = 'b0;
        10'd102 :data = 'b1;
        10'd103 :data = 'b0;
        10'd104 :data = 'b0;
        10'd105 :data = 'b1;
        10'd106 :data = 'b1;
        10'd107 :data = 'b1;
        10'd108 :data = 'b1;
        10'd109 :data = 'b1;
        10'd110 :data = 'b1;
        10'd111 :data = 'b0;
        10'd112 :data = 'b1;
        10'd113 :data = 'b0;
        10'd114 :data = 'b0;
        10'd115 :data = 'b1;
        10'd116 :data = 'b1;
        10'd117 :data = 'b1;
        10'd118 :data = 'b1;
        10'd119 :data = 'b0;
        10'd120 :data = 'b1;
        10'd121 :data = 'b1;
        10'd122 :data = 'b0;
        10'd123 :data = 'b1;
        10'd124 :data = 'b1;
        10'd125 :data = 'b1;
        10'd126 :data = 'b0;
        10'd127 :data = 'b0;
        10'd128 :data = 'b0;
        10'd129 :data = 'b0;
        10'd130 :data = 'b0;
        10'd131 :data = 'b0;
        10'd132 :data = 'b1;
        10'd133 :data = 'b1;
        10'd134 :data = 'b1;
        10'd135 :data = 'b0;
        10'd136 :data = 'b0;
        10'd137 :data = 'b1;
        10'd138 :data = 'b1;
        10'd139 :data = 'b0;
        10'd140 :data = 'b0;
        10'd141 :data = 'b1;
        10'd142 :data = 'b0;
        10'd143 :data = 'b0;
        10'd144 :data = 'b0;
        10'd145 :data = 'b1;
        10'd146 :data = 'b0;
        10'd147 :data = 'b1;
        10'd148 :data = 'b0;
        10'd149 :data = 'b0;
        10'd150 :data = 'b1;
        10'd151 :data = 'b1;
        10'd152 :data = 'b0;
        10'd153 :data = 'b0;
        10'd154 :data = 'b0;
        10'd155 :data = 'b1;
        10'd156 :data = 'b1;
        10'd157 :data = 'b1;
        10'd158 :data = 'b0;
        10'd159 :data = 'b1;
        10'd160 :data = 'b0;
        10'd161 :data = 'b0;
        10'd162 :data = 'b0;
        10'd163 :data = 'b0;
        10'd164 :data = 'b1;
        10'd165 :data = 'b1;
        10'd166 :data = 'b1;
        10'd167 :data = 'b1;
        10'd168 :data = 'b0;
        10'd169 :data = 'b1;
        10'd170 :data = 'b1;
        10'd171 :data = 'b0;
        10'd172 :data = 'b1;
        10'd173 :data = 'b1;
        10'd174 :data = 'b1;
        10'd175 :data = 'b0;
        10'd176 :data = 'b1;
        10'd177 :data = 'b1;
        10'd178 :data = 'b1;
        10'd179 :data = 'b0;
        10'd180 :data = 'b0;
        10'd181 :data = 'b0;
        10'd182 :data = 'b1;
        10'd183 :data = 'b0;
        10'd184 :data = 'b0;
        10'd185 :data = 'b1;
        10'd186 :data = 'b0;
        10'd187 :data = 'b1;
        10'd188 :data = 'b0;
        10'd189 :data = 'b0;
        10'd190 :data = 'b1;
        10'd191 :data = 'b1;
        10'd192 :data = 'b0;
        10'd193 :data = 'b0;
        10'd194 :data = 'b1;
        10'd195 :data = 'b0;
        10'd196 :data = 'b0;
        10'd197 :data = 'b0;
        10'd198 :data = 'b0;
        10'd199 :data = 'b1;
        10'd200 :data = 'b1;
        10'd201 :data = 'b0;
        10'd202 :data = 'b0;
        10'd203 :data = 'b1;
        10'd204 :data = 'b0;
        10'd205 :data = 'b0;
        10'd206 :data = 'b1;
        10'd207 :data = 'b0;
        10'd208 :data = 'b1;
        10'd209 :data = 'b0;
        10'd210 :data = 'b1;
        10'd211 :data = 'b0;
        10'd212 :data = 'b1;
        10'd213 :data = 'b1;
        10'd214 :data = 'b0;
        10'd215 :data = 'b1;
        10'd216 :data = 'b0;
        10'd217 :data = 'b1;
        10'd218 :data = 'b0;
        10'd219 :data = 'b0;
        10'd220 :data = 'b0;
        10'd221 :data = 'b0;
        10'd222 :data = 'b0;
        10'd223 :data = 'b1;
        10'd224 :data = 'b0;
        10'd225 :data = 'b0;
        10'd226 :data = 'b1;
        10'd227 :data = 'b0;
        10'd228 :data = 'b1;
        10'd229 :data = 'b1;
        10'd230 :data = 'b0;
        10'd231 :data = 'b0;
        10'd232 :data = 'b0;
        10'd233 :data = 'b0;
        10'd234 :data = 'b0;
        10'd235 :data = 'b0;
        10'd236 :data = 'b0;
        10'd237 :data = 'b0;
        10'd238 :data = 'b1;
        10'd239 :data = 'b1;
        10'd240 :data = 'b1;
        10'd241 :data = 'b1;
        10'd242 :data = 'b0;
        10'd243 :data = 'b0;
        10'd244 :data = 'b0;
        10'd245 :data = 'b1;
        10'd246 :data = 'b1;
        10'd247 :data = 'b1;
        10'd248 :data = 'b0;
        10'd249 :data = 'b1;
        10'd250 :data = 'b0;
        10'd251 :data = 'b1;
        10'd252 :data = 'b1;
        10'd253 :data = 'b1;
        10'd254 :data = 'b0;
        10'd255 :data = 'b0;
        10'd256 :data = 'b0;
        10'd257 :data = 'b0;
        10'd258 :data = 'b0;
        10'd259 :data = 'b0;
        10'd260 :data = 'b1;
        10'd261 :data = 'b1;
        10'd262 :data = 'b1;
        10'd263 :data = 'b0;
        10'd264 :data = 'b1;
        10'd265 :data = 'b0;
        10'd266 :data = 'b1;
        10'd267 :data = 'b0;
        10'd268 :data = 'b0;
        10'd269 :data = 'b1;
        10'd270 :data = 'b1;
        10'd271 :data = 'b0;
        10'd272 :data = 'b0;
        10'd273 :data = 'b1;
        10'd274 :data = 'b0;
        10'd275 :data = 'b0;
        10'd276 :data = 'b1;
        10'd277 :data = 'b1;
        10'd278 :data = 'b1;
        10'd279 :data = 'b0;
        10'd280 :data = 'b1;
        10'd281 :data = 'b1;
        10'd282 :data = 'b1;
        10'd283 :data = 'b1;
        10'd284 :data = 'b1;
        10'd285 :data = 'b0;
        10'd286 :data = 'b0;
        10'd287 :data = 'b0;
        10'd288 :data = 'b0;
        10'd289 :data = 'b1;
        10'd290 :data = 'b1;
        10'd291 :data = 'b0;
        10'd292 :data = 'b0;
        10'd293 :data = 'b0;
        10'd294 :data = 'b1;
        10'd295 :data = 'b0;
        10'd296 :data = 'b1;
        10'd297 :data = 'b1;
        10'd298 :data = 'b0;
        10'd299 :data = 'b0;
        10'd300 :data = 'b0;
        10'd301 :data = 'b1;
        10'd302 :data = 'b0;
        10'd303 :data = 'b1;
        10'd304 :data = 'b0;
        10'd305 :data = 'b1;
        10'd306 :data = 'b0;
        10'd307 :data = 'b1;
        10'd308 :data = 'b1;
        10'd309 :data = 'b0;
        10'd310 :data = 'b0;
        10'd311 :data = 'b1;
        10'd312 :data = 'b1;
        10'd313 :data = 'b0;
        10'd314 :data = 'b0;
        10'd315 :data = 'b0;
        10'd316 :data = 'b1;
        10'd317 :data = 'b0;
        10'd318 :data = 'b0;
        10'd319 :data = 'b1;
        10'd320 :data = 'b0;
        10'd321 :data = 'b0;
        10'd322 :data = 'b1;
        10'd323 :data = 'b0;
        10'd324 :data = 'b1;
        10'd325 :data = 'b0;
        10'd326 :data = 'b1;
        10'd327 :data = 'b0;
        10'd328 :data = 'b0;
        10'd329 :data = 'b0;
        10'd330 :data = 'b1;
        10'd331 :data = 'b0;
        10'd332 :data = 'b1;
        10'd333 :data = 'b0;
        10'd334 :data = 'b0;
        10'd335 :data = 'b1;
        10'd336 :data = 'b1;
        10'd337 :data = 'b0;
        10'd338 :data = 'b0;
        10'd339 :data = 'b1;
        10'd340 :data = 'b0;
        10'd341 :data = 'b0;
        10'd342 :data = 'b0;
        10'd343 :data = 'b0;
        10'd344 :data = 'b0;
        10'd345 :data = 'b0;
        10'd346 :data = 'b0;
        10'd347 :data = 'b0;
        10'd348 :data = 'b0;
        10'd349 :data = 'b1;
        10'd350 :data = 'b0;
        10'd351 :data = 'b1;
        10'd352 :data = 'b0;
        10'd353 :data = 'b1;
        10'd354 :data = 'b1;
        10'd355 :data = 'b0;
        10'd356 :data = 'b1;
        10'd357 :data = 'b0;
        10'd358 :data = 'b1;
        10'd359 :data = 'b0;
        10'd360 :data = 'b1;
        10'd361 :data = 'b0;
        10'd362 :data = 'b0;
        10'd363 :data = 'b1;
        10'd364 :data = 'b1;
        10'd365 :data = 'b1;
        10'd366 :data = 'b1;
        10'd367 :data = 'b0;
        10'd368 :data = 'b0;
        10'd369 :data = 'b1;
        10'd370 :data = 'b1;
        10'd371 :data = 'b0;
        10'd372 :data = 'b0;
        10'd373 :data = 'b0;
        10'd374 :data = 'b1;
        10'd375 :data = 'b1;
        10'd376 :data = 'b0;
        10'd377 :data = 'b1;
        10'd378 :data = 'b0;
        10'd379 :data = 'b0;
        10'd380 :data = 'b1;
        10'd381 :data = 'b1;
        10'd382 :data = 'b1;
        10'd383 :data = 'b0;
        10'd384 :data = 'b1;
        10'd385 :data = 'b1;
        10'd386 :data = 'b0;
        10'd387 :data = 'b1;
        10'd388 :data = 'b0;
        10'd389 :data = 'b1;
        10'd390 :data = 'b1;
        10'd391 :data = 'b1;
        10'd392 :data = 'b1;
        10'd393 :data = 'b0;
        10'd394 :data = 'b0;
        10'd395 :data = 'b1;
        10'd396 :data = 'b1;
        10'd397 :data = 'b0;
        10'd398 :data = 'b0;
        10'd399 :data = 'b1;
        10'd400 :data = 'b1;
        10'd401 :data = 'b0;
        10'd402 :data = 'b0;
        10'd403 :data = 'b0;
        10'd404 :data = 'b0;
        10'd405 :data = 'b1;
        10'd406 :data = 'b1;
        10'd407 :data = 'b0;
        10'd408 :data = 'b0;
        10'd409 :data = 'b0;
        10'd410 :data = 'b0;
        10'd411 :data = 'b1;
        10'd412 :data = 'b1;
        10'd413 :data = 'b1;
        10'd414 :data = 'b1;
        10'd415 :data = 'b1;
        10'd416 :data = 'b0;
        10'd417 :data = 'b1;
        10'd418 :data = 'b1;
        10'd419 :data = 'b0;
        10'd420 :data = 'b1;
        10'd421 :data = 'b1;
        10'd422 :data = 'b1;
        10'd423 :data = 'b1;
        10'd424 :data = 'b0;
        10'd425 :data = 'b1;
        10'd426 :data = 'b0;
        10'd427 :data = 'b0;
        10'd428 :data = 'b0;
        10'd429 :data = 'b0;
        10'd430 :data = 'b1;
        10'd431 :data = 'b1;
        10'd432 :data = 'b1;
        10'd433 :data = 'b1;
        10'd434 :data = 'b1;
        10'd435 :data = 'b0;
        10'd436 :data = 'b0;
        10'd437 :data = 'b0;
        10'd438 :data = 'b0;
        10'd439 :data = 'b1;
        10'd440 :data = 'b1;
        10'd441 :data = 'b0;
        10'd442 :data = 'b1;
        10'd443 :data = 'b1;
        10'd444 :data = 'b0;
        10'd445 :data = 'b1;
        10'd446 :data = 'b0;
        10'd447 :data = 'b0;
        10'd448 :data = 'b1;
        10'd449 :data = 'b0;
        10'd450 :data = 'b0;
        10'd451 :data = 'b0;
        10'd452 :data = 'b0;
        10'd453 :data = 'b1;
        10'd454 :data = 'b0;
        10'd455 :data = 'b0;
        10'd456 :data = 'b1;
        10'd457 :data = 'b1;
        10'd458 :data = 'b0;
        10'd459 :data = 'b1;
        10'd460 :data = 'b1;
        10'd461 :data = 'b0;
        10'd462 :data = 'b1;
        10'd463 :data = 'b0;
        10'd464 :data = 'b1;
        10'd465 :data = 'b0;
        10'd466 :data = 'b0;
        10'd467 :data = 'b1;
        10'd468 :data = 'b0;
        10'd469 :data = 'b0;
        10'd470 :data = 'b1;
        10'd471 :data = 'b1;
        10'd472 :data = 'b1;
        10'd473 :data = 'b0;
        10'd474 :data = 'b0;
        10'd475 :data = 'b1;
        10'd476 :data = 'b1;
        10'd477 :data = 'b0;
        10'd478 :data = 'b1;
        10'd479 :data = 'b1;
        10'd480 :data = 'b1;
        10'd481 :data = 'b0;
        10'd482 :data = 'b1;
        10'd483 :data = 'b0;
        10'd484 :data = 'b1;
        10'd485 :data = 'b0;
        10'd486 :data = 'b1;
        10'd487 :data = 'b0;
        10'd488 :data = 'b1;
        10'd489 :data = 'b1;
        10'd490 :data = 'b0;
        10'd491 :data = 'b1;
        10'd492 :data = 'b1;
        10'd493 :data = 'b1;
        10'd494 :data = 'b1;
        10'd495 :data = 'b1;
        10'd496 :data = 'b1;
        10'd497 :data = 'b1;
        10'd498 :data = 'b0;
        10'd499 :data = 'b1;
        10'd500 :data = 'b0;
        10'd501 :data = 'b0;
        10'd502 :data = 'b1;
        10'd503 :data = 'b1;
        10'd504 :data = 'b0;
        10'd505 :data = 'b0;
        10'd506 :data = 'b0;
        10'd507 :data = 'b0;
        10'd508 :data = 'b1;
        10'd509 :data = 'b0;
        10'd510 :data = 'b0;
        10'd511 :data = 'b0;
        10'd512 :data = 'b0;
        10'd513 :data = 'b0;
        10'd514 :data = 'b1;
        10'd515 :data = 'b0;
        10'd516 :data = 'b1;
        10'd517 :data = 'b1;
        10'd518 :data = 'b1;
        10'd519 :data = 'b1;
        10'd520 :data = 'b0;
        10'd521 :data = 'b0;
        10'd522 :data = 'b1;
        10'd523 :data = 'b1;
        10'd524 :data = 'b1;
        10'd525 :data = 'b0;
        10'd526 :data = 'b0;
        10'd527 :data = 'b0;
        10'd528 :data = 'b1;
        10'd529 :data = 'b1;
        10'd530 :data = 'b1;
        10'd531 :data = 'b0;
        10'd532 :data = 'b1;
        10'd533 :data = 'b1;
        10'd534 :data = 'b1;
        10'd535 :data = 'b0;
        10'd536 :data = 'b1;
        10'd537 :data = 'b0;
        10'd538 :data = 'b0;
        10'd539 :data = 'b1;
        10'd540 :data = 'b1;
        10'd541 :data = 'b1;
        10'd542 :data = 'b0;
        10'd543 :data = 'b0;
        10'd544 :data = 'b0;
        10'd545 :data = 'b0;
        10'd546 :data = 'b1;
        10'd547 :data = 'b1;
        10'd548 :data = 'b1;
        10'd549 :data = 'b0;
        10'd550 :data = 'b0;
        10'd551 :data = 'b0;
        10'd552 :data = 'b0;
        10'd553 :data = 'b1;
        10'd554 :data = 'b1;
        10'd555 :data = 'b0;
        10'd556 :data = 'b1;
        10'd557 :data = 'b0;
        10'd558 :data = 'b0;
        10'd559 :data = 'b1;
        10'd560 :data = 'b0;
        10'd561 :data = 'b0;
        10'd562 :data = 'b0;
        10'd563 :data = 'b1;
        10'd564 :data = 'b0;
        10'd565 :data = 'b1;
        10'd566 :data = 'b0;
        10'd567 :data = 'b1;
        10'd568 :data = 'b1;
        10'd569 :data = 'b0;
        10'd570 :data = 'b1;
        10'd571 :data = 'b0;
        10'd572 :data = 'b1;
        10'd573 :data = 'b1;
        10'd574 :data = 'b0;
        10'd575 :data = 'b1;
        10'd576 :data = 'b1;
        10'd577 :data = 'b0;
        10'd578 :data = 'b1;
        10'd579 :data = 'b0;
        10'd580 :data = 'b0;
        10'd581 :data = 'b0;
        10'd582 :data = 'b1;
        10'd583 :data = 'b0;
        10'd584 :data = 'b1;
        10'd585 :data = 'b1;
        10'd586 :data = 'b1;
        10'd587 :data = 'b0;
        10'd588 :data = 'b0;
        10'd589 :data = 'b1;
        10'd590 :data = 'b1;
        10'd591 :data = 'b0;
        10'd592 :data = 'b0;
        10'd593 :data = 'b1;
        10'd594 :data = 'b1;
        10'd595 :data = 'b0;
        10'd596 :data = 'b1;
        10'd597 :data = 'b0;
        10'd598 :data = 'b1;
        10'd599 :data = 'b0;
        10'd600 :data = 'b0;
        10'd601 :data = 'b1;
        10'd602 :data = 'b1;
        10'd603 :data = 'b0;
        10'd604 :data = 'b1;
        10'd605 :data = 'b1;
        10'd606 :data = 'b1;
        10'd607 :data = 'b1;
        10'd608 :data = 'b0;
        10'd609 :data = 'b0;
        10'd610 :data = 'b1;
        10'd611 :data = 'b0;
        10'd612 :data = 'b0;
        10'd613 :data = 'b1;
        10'd614 :data = 'b1;
        10'd615 :data = 'b0;
        10'd616 :data = 'b1;
        10'd617 :data = 'b0;
        10'd618 :data = 'b0;
        10'd619 :data = 'b1;
        10'd620 :data = 'b0;
        10'd621 :data = 'b0;
        10'd622 :data = 'b1;
        10'd623 :data = 'b1;
        10'd624 :data = 'b1;
        10'd625 :data = 'b0;
        10'd626 :data = 'b1;
        10'd627 :data = 'b1;
        10'd628 :data = 'b1;
        10'd629 :data = 'b1;
        10'd630 :data = 'b1;
        10'd631 :data = 'b1;
        10'd632 :data = 'b0;
        10'd633 :data = 'b0;
        10'd634 :data = 'b1;
        10'd635 :data = 'b1;
        10'd636 :data = 'b0;
        10'd637 :data = 'b1;
        10'd638 :data = 'b1;
        10'd639 :data = 'b1;
        10'd640 :data = 'b0;
        10'd641 :data = 'b0;
        10'd642 :data = 'b0;
        10'd643 :data = 'b1;
        10'd644 :data = 'b1;
        10'd645 :data = 'b0;
        10'd646 :data = 'b1;
        10'd647 :data = 'b1;
        10'd648 :data = 'b0;
        10'd649 :data = 'b1;
        10'd650 :data = 'b0;
        10'd651 :data = 'b0;
        10'd652 :data = 'b0;
        10'd653 :data = 'b0;
        10'd654 :data = 'b0;
        10'd655 :data = 'b0;
        10'd656 :data = 'b1;
        10'd657 :data = 'b1;
        10'd658 :data = 'b1;
        10'd659 :data = 'b1;
        10'd660 :data = 'b0;
        10'd661 :data = 'b1;
        10'd662 :data = 'b0;
        10'd663 :data = 'b1;
        10'd664 :data = 'b1;
        10'd665 :data = 'b0;
        10'd666 :data = 'b1;
        10'd667 :data = 'b0;
        10'd668 :data = 'b0;
        10'd669 :data = 'b0;
        10'd670 :data = 'b1;
        10'd671 :data = 'b0;
        10'd672 :data = 'b1;
        10'd673 :data = 'b0;
        10'd674 :data = 'b1;
        10'd675 :data = 'b1;
        10'd676 :data = 'b1;
        10'd677 :data = 'b0;
        10'd678 :data = 'b1;
        10'd679 :data = 'b1;
        10'd680 :data = 'b0;
        10'd681 :data = 'b1;
        10'd682 :data = 'b1;
        10'd683 :data = 'b1;
        10'd684 :data = 'b1;
        10'd685 :data = 'b1;
        10'd686 :data = 'b1;
        10'd687 :data = 'b0;
        10'd688 :data = 'b0;
        10'd689 :data = 'b0;
        10'd690 :data = 'b0;
        10'd691 :data = 'b1;
        10'd692 :data = 'b0;
        10'd693 :data = 'b1;
        10'd694 :data = 'b1;
        10'd695 :data = 'b1;
        10'd696 :data = 'b1;
        10'd697 :data = 'b0;
        10'd698 :data = 'b0;
        10'd699 :data = 'b0;
        10'd700 :data = 'b0;
        10'd701 :data = 'b1;
        10'd702 :data = 'b1;
        10'd703 :data = 'b1;
        10'd704 :data = 'b0;
        10'd705 :data = 'b0;
        10'd706 :data = 'b1;
        10'd707 :data = 'b1;
        10'd708 :data = 'b0;
        10'd709 :data = 'b0;
        10'd710 :data = 'b0;
        10'd711 :data = 'b1;
        10'd712 :data = 'b1;
        10'd713 :data = 'b1;
        10'd714 :data = 'b1;
        10'd715 :data = 'b0;
        10'd716 :data = 'b1;
        10'd717 :data = 'b1;
        10'd718 :data = 'b1;
        10'd719 :data = 'b1;
        10'd720 :data = 'b0;
        10'd721 :data = 'b0;
        10'd722 :data = 'b0;
        10'd723 :data = 'b0;
        10'd724 :data = 'b1;
        10'd725 :data = 'b0;
        10'd726 :data = 'b1;
        10'd727 :data = 'b1;
        10'd728 :data = 'b0;
        10'd729 :data = 'b0;
        10'd730 :data = 'b0;
        10'd731 :data = 'b1;
        10'd732 :data = 'b1;
        10'd733 :data = 'b1;
        10'd734 :data = 'b0;
        10'd735 :data = 'b0;
        10'd736 :data = 'b0;
        10'd737 :data = 'b1;
        10'd738 :data = 'b1;
        10'd739 :data = 'b0;
        10'd740 :data = 'b1;
        10'd741 :data = 'b0;
        10'd742 :data = 'b0;
        10'd743 :data = 'b1;
        10'd744 :data = 'b1;
        10'd745 :data = 'b0;
        10'd746 :data = 'b0;
        10'd747 :data = 'b0;
        10'd748 :data = 'b1;
        10'd749 :data = 'b0;
        10'd750 :data = 'b0;
        10'd751 :data = 'b0;
        10'd752 :data = 'b0;
        10'd753 :data = 'b1;
        10'd754 :data = 'b0;
        10'd755 :data = 'b0;
        10'd756 :data = 'b1;
        10'd757 :data = 'b1;
        10'd758 :data = 'b0;
        10'd759 :data = 'b0;
        10'd760 :data = 'b1;
        10'd761 :data = 'b0;
        10'd762 :data = 'b1;
        10'd763 :data = 'b1;
        10'd764 :data = 'b1;
        10'd765 :data = 'b1;
        10'd766 :data = 'b1;
        10'd767 :data = 'b0;
        10'd768 :data = 'b0;
        10'd769 :data = 'b1;
        10'd770 :data = 'b1;
        10'd771 :data = 'b0;
        10'd772 :data = 'b1;
        10'd773 :data = 'b0;
        10'd774 :data = 'b0;
        10'd775 :data = 'b1;
        10'd776 :data = 'b1;
        10'd777 :data = 'b1;
        10'd778 :data = 'b0;
        10'd779 :data = 'b0;
        10'd780 :data = 'b0;
        10'd781 :data = 'b1;
        10'd782 :data = 'b0;
        10'd783 :data = 'b0;
        10'd784 :data = 'b0;
        10'd785 :data = 'b0;
        10'd786 :data = 'b1;
        10'd787 :data = 'b1;
        10'd788 :data = 'b1;
        10'd789 :data = 'b0;
        10'd790 :data = 'b1;
        10'd791 :data = 'b1;
        10'd792 :data = 'b1;
        10'd793 :data = 'b0;
        10'd794 :data = 'b0;
        10'd795 :data = 'b1;
        10'd796 :data = 'b1;
        10'd797 :data = 'b0;
        10'd798 :data = 'b1;
        10'd799 :data = 'b0;
        10'd800 :data = 'b0;
        10'd801 :data = 'b1;
        10'd802 :data = 'b1;
        10'd803 :data = 'b0;
        10'd804 :data = 'b0;
        10'd805 :data = 'b0;
        10'd806 :data = 'b1;
        10'd807 :data = 'b0;
        10'd808 :data = 'b0;
        10'd809 :data = 'b1;
        10'd810 :data = 'b0;
        10'd811 :data = 'b0;
        10'd812 :data = 'b1;
        10'd813 :data = 'b1;
        10'd814 :data = 'b0;
        10'd815 :data = 'b1;
        10'd816 :data = 'b0;
        10'd817 :data = 'b0;
        10'd818 :data = 'b0;
        10'd819 :data = 'b1;
        10'd820 :data = 'b0;
        10'd821 :data = 'b0;
        10'd822 :data = 'b1;
        10'd823 :data = 'b1;
        10'd824 :data = 'b0;
        10'd825 :data = 'b1;
        10'd826 :data = 'b1;
        10'd827 :data = 'b0;
        10'd828 :data = 'b1;
        10'd829 :data = 'b0;
        10'd830 :data = 'b0;
        10'd831 :data = 'b0;
        10'd832 :data = 'b0;
        10'd833 :data = 'b0;
        10'd834 :data = 'b0;
        10'd835 :data = 'b1;
        10'd836 :data = 'b0;
        10'd837 :data = 'b1;
        10'd838 :data = 'b1;
        10'd839 :data = 'b1;
        10'd840 :data = 'b0;
        10'd841 :data = 'b1;
        10'd842 :data = 'b0;
        10'd843 :data = 'b1;
        10'd844 :data = 'b0;
        10'd845 :data = 'b1;
        10'd846 :data = 'b0;
        10'd847 :data = 'b1;
        10'd848 :data = 'b1;
        10'd849 :data = 'b0;
        10'd850 :data = 'b0;
        10'd851 :data = 'b0;
        10'd852 :data = 'b1;
        10'd853 :data = 'b0;
        10'd854 :data = 'b1;
        10'd855 :data = 'b0;
        10'd856 :data = 'b0;
        10'd857 :data = 'b1;
        10'd858 :data = 'b1;
        10'd859 :data = 'b1;
        10'd860 :data = 'b0;
        10'd861 :data = 'b0;
        10'd862 :data = 'b1;
        10'd863 :data = 'b1;
        10'd864 :data = 'b1;
        10'd865 :data = 'b1;
        10'd866 :data = 'b0;
        10'd867 :data = 'b0;
        10'd868 :data = 'b0;
        10'd869 :data = 'b1;
        10'd870 :data = 'b1;
        10'd871 :data = 'b0;
        10'd872 :data = 'b0;
        10'd873 :data = 'b1;
        10'd874 :data = 'b0;
        10'd875 :data = 'b1;
        10'd876 :data = 'b1;
        10'd877 :data = 'b0;
        10'd878 :data = 'b1;
        10'd879 :data = 'b0;
        10'd880 :data = 'b1;
        10'd881 :data = 'b0;
        10'd882 :data = 'b0;
        10'd883 :data = 'b0;
        10'd884 :data = 'b1;
        10'd885 :data = 'b1;
        10'd886 :data = 'b0;
        10'd887 :data = 'b1;
        10'd888 :data = 'b0;
        10'd889 :data = 'b1;
        10'd890 :data = 'b1;
        10'd891 :data = 'b1;
        10'd892 :data = 'b1;
        10'd893 :data = 'b0;
        10'd894 :data = 'b0;
        10'd895 :data = 'b1;
        10'd896 :data = 'b1;
        10'd897 :data = 'b0;
        10'd898 :data = 'b1;
        10'd899 :data = 'b0;
        10'd900 :data = 'b0;
        10'd901 :data = 'b1;
        10'd902 :data = 'b0;
        10'd903 :data = 'b1;
        10'd904 :data = 'b0;
        10'd905 :data = 'b1;
        10'd906 :data = 'b0;
        10'd907 :data = 'b0;
        10'd908 :data = 'b0;
        10'd909 :data = 'b1;
        10'd910 :data = 'b1;
        10'd911 :data = 'b0;
        10'd912 :data = 'b1;
        10'd913 :data = 'b1;
        10'd914 :data = 'b0;
        10'd915 :data = 'b0;
        10'd916 :data = 'b1;
        10'd917 :data = 'b0;
        10'd918 :data = 'b1;
        10'd919 :data = 'b0;
        10'd920 :data = 'b1;
        10'd921 :data = 'b1;
        10'd922 :data = 'b0;
        10'd923 :data = 'b1;
        10'd924 :data = 'b0;
        10'd925 :data = 'b1;
        10'd926 :data = 'b1;
        10'd927 :data = 'b1;
        10'd928 :data = 'b1;
        10'd929 :data = 'b1;
        10'd930 :data = 'b0;
        10'd931 :data = 'b0;
        10'd932 :data = 'b0;
        10'd933 :data = 'b0;
        10'd934 :data = 'b0;
        10'd935 :data = 'b1;
        10'd936 :data = 'b1;
        10'd937 :data = 'b1;
        10'd938 :data = 'b0;
        10'd939 :data = 'b1;
        10'd940 :data = 'b1;
        10'd941 :data = 'b1;
        10'd942 :data = 'b0;
        10'd943 :data = 'b0;
        10'd944 :data = 'b0;
        10'd945 :data = 'b0;
        10'd946 :data = 'b1;
        10'd947 :data = 'b1;
        10'd948 :data = 'b0;
        10'd949 :data = 'b0;
        10'd950 :data = 'b0;
        10'd951 :data = 'b1;
        10'd952 :data = 'b0;
        10'd953 :data = 'b1;
        10'd954 :data = 'b1;
        10'd955 :data = 'b1;
        10'd956 :data = 'b1;
        10'd957 :data = 'b0;
        10'd958 :data = 'b1;
        10'd959 :data = 'b1;
        10'd960 :data = 'b1;
        10'd961 :data = 'b0;
        10'd962 :data = 'b0;
        10'd963 :data = 'b1;
        10'd964 :data = 'b0;
        10'd965 :data = 'b1;
        10'd966 :data = 'b1;
        10'd967 :data = 'b1;
        10'd968 :data = 'b0;
        10'd969 :data = 'b1;
        10'd970 :data = 'b0;
        10'd971 :data = 'b0;
        10'd972 :data = 'b1;
        10'd973 :data = 'b0;
        10'd974 :data = 'b0;
        10'd975 :data = 'b0;
        10'd976 :data = 'b1;
        10'd977 :data = 'b1;
        10'd978 :data = 'b0;
        10'd979 :data = 'b0;
        10'd980 :data = 'b0;
        10'd981 :data = 'b1;
        10'd982 :data = 'b1;
        10'd983 :data = 'b1;
        10'd984 :data = 'b1;
        10'd985 :data = 'b0;
        10'd986 :data = 'b0;
        10'd987 :data = 'b0;
        10'd988 :data = 'b1;
        10'd989 :data = 'b0;
        10'd990 :data = 'b0;
        10'd991 :data = 'b0;
        10'd992 :data = 'b0;
        10'd993 :data = 'b1;
        10'd994 :data = 'b1;
        10'd995 :data = 'b0;
        10'd996 :data = 'b1;
        10'd997 :data = 'b1;
        10'd998 :data = 'b0;
        10'd999 :data = 'b0;
        10'd1000 :data = 'b1;
        10'd1001 :data = 'b1;
        10'd1002 :data = 'b1;
        10'd1003 :data = 'b1;
        10'd1004 :data = 'b1;
        10'd1005 :data = 'b1;
        10'd1006 :data = 'b0;
        10'd1007 :data = 'b1;
        10'd1008 :data = 'b1;
        10'd1009 :data = 'b1;
        10'd1010 :data = 'b0;
        10'd1011 :data = 'b1;
        10'd1012 :data = 'b1;
        10'd1013 :data = 'b1;
        10'd1014 :data = 'b0;
        10'd1015 :data = 'b0;
        10'd1016 :data = 'b1;
        10'd1017 :data = 'b1;
        10'd1018 :data = 'b1;
        10'd1019 :data = 'b1;
        10'd1020 :data = 'b1;
        10'd1021 :data = 'b1;
        10'd1022 :data = 'b0;
        10'd1023 :data = 'b0;
        default: data = 'b0;
    endcase
end

endmodule
